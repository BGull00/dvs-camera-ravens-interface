`ifndef DVS_RAVENS_PKG
    `define DVS_RAVENS_PKG

    package dvs_ravens_pkg;

        localparam DVS_WIDTH_PXLS = 346;
        localparam DVS_HEIGHT_PXLS = 260;

    endpackage: dvs_ravens_pkg