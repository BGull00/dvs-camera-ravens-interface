module sram_compiled_array(addr0,addr1,addr2,addr3,addr4,addr5,addr6,addr7,addr8,addr9,din0,din1,din2,din3,din4,din5,din6,din7,din8,din9,din10,din11,din12,din13,din14,din15,din16,din17,din18,din19,din20,din21,din22,din23,din24,din25,din26,din27,din28,din29,din30,din31,din32,din33,din34,din35,din36,din37,din38,din39,din40,din41,din42,din43,din44,din45,din46,din47,din48,din49,din50,din51,din52,din53,din54,din55,din56,din57,din58,din59,din60,din61,din62,din63,dout0,dout1,dout2,dout3,dout4,dout5,dout6,dout7,dout8,dout9,dout10,dout11,dout12,dout13,dout14,dout15,dout16,dout17,dout18,dout19,dout20,dout21,dout22,dout23,dout24,dout25,dout26,dout27,dout28,dout29,dout30,dout31,dout32,dout33,dout34,dout35,dout36,dout37,dout38,dout39,dout40,dout41,dout42,dout43,dout44,dout45,dout46,dout47,dout48,dout49,dout50,dout51,dout52,dout53,dout54,dout55,dout56,dout57,dout58,dout59,dout60,dout61,dout62,dout63,clk,write_en,sense_en);
endmodule: sram_compiled_array