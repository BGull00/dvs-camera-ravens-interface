module sram_compiled_array(addr0,addr1,addr2,addr3,addr4,addr5,addr6,addr7,addr8,addr9,din0,din1,din2,din3,din4,din5,din6,din7,din8,din9,din10,din11,din12,din13,din14,din15,din16,din17,din18,din19,din20,din21,din22,din23,din24,din25,din26,din27,din28,din29,din30,din31,din32,din33,din34,din35,din36,din37,din38,din39,din40,din41,din42,din43,din44,din45,din46,din47,din48,din49,din50,din51,din52,din53,din54,din55,din56,din57,din58,din59,din60,din61,din62,din63,dout0,dout1,dout2,dout3,dout4,dout5,dout6,dout7,dout8,dout9,dout10,dout11,dout12,dout13,dout14,dout15,dout16,dout17,dout18,dout19,dout20,dout21,dout22,dout23,dout24,dout25,dout26,dout27,dout28,dout29,dout30,dout31,dout32,dout33,dout34,dout35,dout36,dout37,dout38,dout39,dout40,dout41,dout42,dout43,dout44,dout45,dout46,dout47,dout48,dout49,dout50,dout51,dout52,dout53,dout54,dout55,dout56,dout57,dout58,dout59,dout60,dout61,dout62,dout63,clk,write_en,sense_en);
    input addr0;
    input addr1;
    input addr2;
    input addr3;
    input addr4;
    input addr5;
    input addr6;
    input addr7;
    input addr8;
    input addr9;
    input din0;
    input din1;
    input din2;
    input din3;
    input din4;
    input din5;
    input din6;
    input din7;
    input din8;
    input din9;
    input din10;
    input din11;
    input din12;
    input din13;
    input din14;
    input din15;
    input din16;
    input din17;
    input din18;
    input din19;
    input din20;
    input din21;
    input din22;
    input din23;
    input din24;
    input din25;
    input din26;
    input din27;
    input din28;
    input din29;
    input din30;
    input din31;
    input din32;
    input din33;
    input din34;
    input din35;
    input din36;
    input din37;
    input din38;
    input din39;
    input din40;
    input din41;
    input din42;
    input din43;
    input din44;
    input din45;
    input din46;
    input din47;
    input din48;
    input din49;
    input din50;
    input din51;
    input din52;
    input din53;
    input din54;
    input din55;
    input din56;
    input din57;
    input din58;
    input din59;
    input din60;
    input din61;
    input din62;
    input din63;
    output dout0;
    output dout1;
    output dout2;
    output dout3;
    output dout4;
    output dout5;
    output dout6;
    output dout7;
    output dout8;
    output dout9;
    output dout10;
    output dout11;
    output dout12;
    output dout13;
    output dout14;
    output dout15;
    output dout16;
    output dout17;
    output dout18;
    output dout19;
    output dout20;
    output dout21;
    output dout22;
    output dout23;
    output dout24;
    output dout25;
    output dout26;
    output dout27;
    output dout28;
    output dout29;
    output dout30;
    output dout31;
    output dout32;
    output dout33;
    output dout34;
    output dout35;
    output dout36;
    output dout37;
    output dout38;
    output dout39;
    output dout40;
    output dout41;
    output dout42;
    output dout43;
    output dout44;
    output dout45;
    output dout46;
    output dout47;
    output dout48;
    output dout49;
    output dout50;
    output dout51;
    output dout52;
    output dout53;
    output dout54;
    output dout55;
    output dout56;
    output dout57;
    output dout58;
    output dout59;
    output dout60;
    output dout61;
    output dout62;
    output dout63;
    input clk;
    input write_en;
    input sense_en;
endmodule: sram_compiled_array