VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_compiled_array
  CLASS CORE ;
  ORIGIN 33.525 68.925 ;
  FOREIGN sram_compiled_array -33.525 -68.925 ;
  SIZE 76.79 BY 78.82 ;
  SYMMETRY X Y ;
  SITE CoreSite ;
  PIN write_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.235 -59.445 36.83 -59.355 ;
        RECT 36.65 -59.535 36.83 -59.355 ;
        RECT 31.85 -59.535 32.03 -59.355 ;
        RECT 27.05 -59.535 27.23 -59.355 ;
        RECT 22.25 -59.535 22.43 -59.355 ;
        RECT 17.45 -59.535 17.63 -59.355 ;
        RECT 12.65 -59.535 12.83 -59.355 ;
        RECT 7.85 -59.535 8.03 -59.355 ;
        RECT 3.05 -59.535 3.23 -59.355 ;
    END
  END write_en
  PIN din0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.29 -59.765 -0.06 -59.535 ;
      LAYER M3 ;
        RECT -0.29 -59.765 -0.06 -59.535 ;
      LAYER M1 ;
        RECT -0.29 -59.625 1.625 -59.535 ;
        RECT -0.29 -59.765 -0.06 -59.535 ;
      LAYER V2 ;
        RECT -0.225 -59.7 -0.125 -59.6 ;
      LAYER V1 ;
        RECT -0.225 -59.7 -0.125 -59.6 ;
    END
  END din0
  PIN din1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 4.51 -59.765 4.74 -59.535 ;
      LAYER M3 ;
        RECT 4.51 -59.765 4.74 -59.535 ;
      LAYER M1 ;
        RECT 4.51 -59.625 6.425 -59.535 ;
        RECT 4.51 -59.765 4.74 -59.535 ;
      LAYER V2 ;
        RECT 4.575 -59.7 4.675 -59.6 ;
      LAYER V1 ;
        RECT 4.575 -59.7 4.675 -59.6 ;
    END
  END din1
  PIN din2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 9.31 -59.765 9.54 -59.535 ;
      LAYER M3 ;
        RECT 9.31 -59.765 9.54 -59.535 ;
      LAYER M1 ;
        RECT 9.31 -59.625 11.225 -59.535 ;
        RECT 9.31 -59.765 9.54 -59.535 ;
      LAYER V2 ;
        RECT 9.375 -59.7 9.475 -59.6 ;
      LAYER V1 ;
        RECT 9.375 -59.7 9.475 -59.6 ;
    END
  END din2
  PIN din3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 14.11 -59.765 14.34 -59.535 ;
      LAYER M3 ;
        RECT 14.11 -59.765 14.34 -59.535 ;
      LAYER M1 ;
        RECT 14.11 -59.625 16.025 -59.535 ;
        RECT 14.11 -59.765 14.34 -59.535 ;
      LAYER V2 ;
        RECT 14.175 -59.7 14.275 -59.6 ;
      LAYER V1 ;
        RECT 14.175 -59.7 14.275 -59.6 ;
    END
  END din3
  PIN din4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.91 -59.765 19.14 -59.535 ;
      LAYER M3 ;
        RECT 18.91 -59.765 19.14 -59.535 ;
      LAYER M1 ;
        RECT 18.91 -59.625 20.825 -59.535 ;
        RECT 18.91 -59.765 19.14 -59.535 ;
      LAYER V2 ;
        RECT 18.975 -59.7 19.075 -59.6 ;
      LAYER V1 ;
        RECT 18.975 -59.7 19.075 -59.6 ;
    END
  END din4
  PIN din5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.71 -59.765 23.94 -59.535 ;
      LAYER M3 ;
        RECT 23.71 -59.765 23.94 -59.535 ;
      LAYER M1 ;
        RECT 23.71 -59.625 25.625 -59.535 ;
        RECT 23.71 -59.765 23.94 -59.535 ;
      LAYER V2 ;
        RECT 23.775 -59.7 23.875 -59.6 ;
      LAYER V1 ;
        RECT 23.775 -59.7 23.875 -59.6 ;
    END
  END din5
  PIN din6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 28.51 -59.765 28.74 -59.535 ;
      LAYER M3 ;
        RECT 28.51 -59.765 28.74 -59.535 ;
      LAYER M1 ;
        RECT 28.51 -59.625 30.425 -59.535 ;
        RECT 28.51 -59.765 28.74 -59.535 ;
      LAYER V2 ;
        RECT 28.575 -59.7 28.675 -59.6 ;
      LAYER V1 ;
        RECT 28.575 -59.7 28.675 -59.6 ;
    END
  END din6
  PIN din7
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.31 -59.765 33.54 -59.535 ;
      LAYER M3 ;
        RECT 33.31 -59.765 33.54 -59.535 ;
      LAYER M1 ;
        RECT 33.31 -59.625 35.225 -59.535 ;
        RECT 33.31 -59.765 33.54 -59.535 ;
      LAYER V2 ;
        RECT 33.375 -59.7 33.475 -59.6 ;
      LAYER V1 ;
        RECT 33.375 -59.7 33.475 -59.6 ;
    END
  END din7
  PIN sense_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -0.03 -62.425 34.535 -62.305 ;
    END
  END sense_en
  PIN dout0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 1.95 -62.17 2.05 -61.42 ;
        RECT -0.03 -62.115 2.05 -61.995 ;
        RECT 1.58 -62.17 2.05 -61.995 ;
        RECT 0.405 -62.115 0.505 -61.41 ;
    END
  END dout0
  PIN dout1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 6.75 -62.17 6.85 -61.42 ;
        RECT 4.77 -62.115 6.85 -61.995 ;
        RECT 6.38 -62.17 6.85 -61.995 ;
        RECT 5.205 -62.115 5.305 -61.41 ;
    END
  END dout1
  PIN dout2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 11.55 -62.17 11.65 -61.42 ;
        RECT 9.57 -62.115 11.65 -61.995 ;
        RECT 11.18 -62.17 11.65 -61.995 ;
        RECT 10.005 -62.115 10.105 -61.41 ;
    END
  END dout2
  PIN dout3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 16.35 -62.17 16.45 -61.42 ;
        RECT 14.37 -62.115 16.45 -61.995 ;
        RECT 15.98 -62.17 16.45 -61.995 ;
        RECT 14.805 -62.115 14.905 -61.41 ;
    END
  END dout3
  PIN dout4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 21.15 -62.17 21.25 -61.42 ;
        RECT 19.17 -62.115 21.25 -61.995 ;
        RECT 20.78 -62.17 21.25 -61.995 ;
        RECT 19.605 -62.115 19.705 -61.41 ;
    END
  END dout4
  PIN dout5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 25.95 -62.17 26.05 -61.42 ;
        RECT 23.97 -62.115 26.05 -61.995 ;
        RECT 25.58 -62.17 26.05 -61.995 ;
        RECT 24.405 -62.115 24.505 -61.41 ;
    END
  END dout5
  PIN dout6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 30.75 -62.17 30.85 -61.42 ;
        RECT 28.77 -62.115 30.85 -61.995 ;
        RECT 30.38 -62.17 30.85 -61.995 ;
        RECT 29.205 -62.115 29.305 -61.41 ;
    END
  END dout6
  PIN dout7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT 35.55 -62.17 35.65 -61.42 ;
        RECT 33.57 -62.115 35.65 -61.995 ;
        RECT 35.18 -62.17 35.65 -61.995 ;
        RECT 34.005 -62.115 34.105 -61.41 ;
    END
  END dout7
  PIN gnd!
    DIRECTION INPUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 42.265 -64.965 43.265 9.895 ;
        RECT 38.4 -50.165 38.5 9.895 ;
        RECT 37.2 -50.165 37.3 9.895 ;
        RECT 36 -50.165 36.1 9.895 ;
        RECT 34.8 -50.165 34.9 9.895 ;
        RECT 33.6 -50.165 33.7 9.895 ;
        RECT 32.4 -50.165 32.5 9.895 ;
        RECT 31.2 -50.165 31.3 9.895 ;
        RECT 30 -50.165 30.1 9.895 ;
        RECT 28.8 -50.165 28.9 9.895 ;
        RECT 27.6 -50.165 27.7 9.895 ;
        RECT 26.4 -50.165 26.5 9.895 ;
        RECT 25.2 -50.165 25.3 9.895 ;
        RECT 24 -50.165 24.1 9.895 ;
        RECT 22.8 -50.165 22.9 9.895 ;
        RECT 21.6 -50.165 21.7 9.895 ;
        RECT 20.4 -50.165 20.5 9.895 ;
        RECT 19.2 -50.165 19.3 9.895 ;
        RECT 18 -50.165 18.1 9.895 ;
        RECT 16.8 -50.165 16.9 9.895 ;
        RECT 15.6 -50.165 15.7 9.895 ;
        RECT 14.4 -50.165 14.5 9.895 ;
        RECT 13.2 -50.165 13.3 9.895 ;
        RECT 12 -50.165 12.1 9.895 ;
        RECT 10.8 -50.165 10.9 9.895 ;
        RECT 9.6 -50.165 9.7 9.895 ;
        RECT 8.4 -50.165 8.5 9.895 ;
        RECT 7.2 -50.165 7.3 9.895 ;
        RECT 6 -50.165 6.1 9.895 ;
        RECT 4.8 -50.165 4.9 9.895 ;
        RECT 3.6 -50.165 3.7 9.895 ;
        RECT 2.4 -50.165 2.5 9.895 ;
        RECT 1.2 -50.165 1.3 9.895 ;
        RECT 0 -50.165 0.1 9.895 ;
        RECT -1.805 -55.975 -1.705 -55.375 ;
        RECT -1.805 -44.755 -1.705 -44.155 ;
        RECT -1.805 -43.055 -1.705 -42.455 ;
        RECT -1.805 -31.835 -1.705 -31.235 ;
        RECT -1.805 -30.135 -1.705 -29.535 ;
        RECT -1.805 -18.915 -1.705 -18.315 ;
        RECT -1.805 -17.215 -1.705 -16.615 ;
        RECT -1.805 -5.995 -1.705 -5.395 ;
        RECT -1.805 -4.295 -1.705 -3.695 ;
        RECT -3.105 -55.975 -3.005 -55.375 ;
        RECT -3.105 -44.755 -3.005 -44.155 ;
        RECT -3.105 -43.055 -3.005 -42.455 ;
        RECT -3.105 -31.835 -3.005 -31.235 ;
        RECT -3.105 -30.135 -3.005 -29.535 ;
        RECT -3.105 -18.915 -3.005 -18.315 ;
        RECT -3.105 -17.215 -3.005 -16.615 ;
        RECT -3.105 -5.995 -3.005 -5.395 ;
        RECT -3.105 -4.295 -3.005 -3.695 ;
        RECT -4.405 -55.975 -4.305 -55.375 ;
        RECT -4.405 -44.755 -4.305 -44.155 ;
        RECT -4.405 -43.055 -4.305 -42.455 ;
        RECT -4.405 -31.835 -4.305 -31.235 ;
        RECT -4.405 -30.135 -4.305 -29.535 ;
        RECT -4.405 -18.915 -4.305 -18.315 ;
        RECT -4.405 -17.215 -4.305 -16.615 ;
        RECT -4.405 -5.995 -4.305 -5.395 ;
        RECT -4.405 -4.295 -4.305 -3.695 ;
        RECT -5.705 -55.975 -5.605 -55.375 ;
        RECT -5.705 -44.755 -5.605 -44.155 ;
        RECT -5.705 -43.055 -5.605 -42.455 ;
        RECT -5.705 -31.835 -5.605 -31.235 ;
        RECT -5.705 -30.135 -5.605 -29.535 ;
        RECT -5.705 -18.915 -5.605 -18.315 ;
        RECT -5.705 -17.215 -5.605 -16.615 ;
        RECT -5.705 -5.995 -5.605 -5.395 ;
        RECT -5.705 -4.295 -5.605 -3.695 ;
        RECT -33.525 -63.475 -32.525 9.895 ;
      LAYER M1 ;
        RECT 6 -6.065 6.1 -5.53 ;
        RECT 6 -4.16 6.1 -3.625 ;
        RECT 6 -2.835 6.1 -2.3 ;
        RECT 6 -0.93 6.1 -0.395 ;
        RECT 6 0.395 6.1 0.93 ;
        RECT 4.8 -49.38 4.9 -48.845 ;
        RECT 4.8 -48.055 4.9 -47.52 ;
        RECT 4.8 -46.15 4.9 -45.615 ;
        RECT 4.8 -44.825 4.9 -44.29 ;
        RECT 4.8 -42.92 4.9 -42.385 ;
        RECT 4.8 -41.595 4.9 -41.06 ;
        RECT 4.8 -39.69 4.9 -39.155 ;
        RECT 4.8 -38.365 4.9 -37.83 ;
        RECT 4.8 -36.46 4.9 -35.925 ;
        RECT 4.8 -35.135 4.9 -34.6 ;
        RECT 4.8 -33.23 4.9 -32.695 ;
        RECT 4.8 -31.905 4.9 -31.37 ;
        RECT 4.8 -30 4.9 -29.465 ;
        RECT 4.8 -28.675 4.9 -28.14 ;
        RECT 4.8 -26.77 4.9 -26.235 ;
        RECT 4.8 -25.445 4.9 -24.91 ;
        RECT 4.8 -23.54 4.9 -23.005 ;
        RECT 4.8 -22.215 4.9 -21.68 ;
        RECT 4.8 -20.31 4.9 -19.775 ;
        RECT 4.8 -18.985 4.9 -18.45 ;
        RECT 4.8 -17.08 4.9 -16.545 ;
        RECT 4.8 -15.755 4.9 -15.22 ;
        RECT 4.8 -13.85 4.9 -13.315 ;
        RECT 4.8 -12.525 4.9 -11.99 ;
        RECT 4.8 -10.62 4.9 -10.085 ;
        RECT 4.8 -9.295 4.9 -8.76 ;
        RECT 4.8 -7.39 4.9 -6.855 ;
        RECT 4.8 -6.065 4.9 -5.53 ;
        RECT 4.8 -4.16 4.9 -3.625 ;
        RECT 4.8 -2.835 4.9 -2.3 ;
        RECT 4.8 -0.93 4.9 -0.395 ;
        RECT 4.8 0.395 4.9 0.93 ;
        RECT 3.6 -49.38 3.7 -48.845 ;
        RECT 3.6 -48.055 3.7 -47.52 ;
        RECT 3.6 -46.15 3.7 -45.615 ;
        RECT 3.6 -44.825 3.7 -44.29 ;
        RECT 3.6 -42.92 3.7 -42.385 ;
        RECT 3.6 -41.595 3.7 -41.06 ;
        RECT 3.6 -39.69 3.7 -39.155 ;
        RECT 3.6 -38.365 3.7 -37.83 ;
        RECT 3.6 -36.46 3.7 -35.925 ;
        RECT 3.6 -35.135 3.7 -34.6 ;
        RECT 3.6 -33.23 3.7 -32.695 ;
        RECT 3.6 -31.905 3.7 -31.37 ;
        RECT 3.6 -30 3.7 -29.465 ;
        RECT 3.6 -28.675 3.7 -28.14 ;
        RECT 3.6 -26.77 3.7 -26.235 ;
        RECT 3.6 -25.445 3.7 -24.91 ;
        RECT 3.6 -23.54 3.7 -23.005 ;
        RECT 3.6 -22.215 3.7 -21.68 ;
        RECT 3.6 -20.31 3.7 -19.775 ;
        RECT 3.6 -18.985 3.7 -18.45 ;
        RECT 3.6 -17.08 3.7 -16.545 ;
        RECT 3.6 -15.755 3.7 -15.22 ;
        RECT 3.6 -13.85 3.7 -13.315 ;
        RECT 3.6 -12.525 3.7 -11.99 ;
        RECT 3.6 -10.62 3.7 -10.085 ;
        RECT 3.6 -9.295 3.7 -8.76 ;
        RECT 3.6 -7.39 3.7 -6.855 ;
        RECT 3.6 -6.065 3.7 -5.53 ;
        RECT 3.6 -4.16 3.7 -3.625 ;
        RECT 3.6 -2.835 3.7 -2.3 ;
        RECT 3.6 -0.93 3.7 -0.395 ;
        RECT 3.6 0.395 3.7 0.93 ;
        RECT 2.4 -49.38 2.5 -48.845 ;
        RECT 2.4 -48.055 2.5 -47.52 ;
        RECT 2.4 -46.15 2.5 -45.615 ;
        RECT 2.4 -44.825 2.5 -44.29 ;
        RECT 2.4 -42.92 2.5 -42.385 ;
        RECT 2.4 -41.595 2.5 -41.06 ;
        RECT 2.4 -39.69 2.5 -39.155 ;
        RECT 2.4 -38.365 2.5 -37.83 ;
        RECT 2.4 -36.46 2.5 -35.925 ;
        RECT 2.4 -35.135 2.5 -34.6 ;
        RECT 2.4 -33.23 2.5 -32.695 ;
        RECT 2.4 -31.905 2.5 -31.37 ;
        RECT 2.4 -30 2.5 -29.465 ;
        RECT 2.4 -28.675 2.5 -28.14 ;
        RECT 2.4 -26.77 2.5 -26.235 ;
        RECT 2.4 -25.445 2.5 -24.91 ;
        RECT 2.4 -23.54 2.5 -23.005 ;
        RECT 2.4 -22.215 2.5 -21.68 ;
        RECT 2.4 -20.31 2.5 -19.775 ;
        RECT 2.4 -18.985 2.5 -18.45 ;
        RECT 2.4 -17.08 2.5 -16.545 ;
        RECT 2.4 -15.755 2.5 -15.22 ;
        RECT 2.4 -13.85 2.5 -13.315 ;
        RECT 2.4 -12.525 2.5 -11.99 ;
        RECT 2.4 -10.62 2.5 -10.085 ;
        RECT 2.4 -9.295 2.5 -8.76 ;
        RECT 2.4 -7.39 2.5 -6.855 ;
        RECT 2.4 -6.065 2.5 -5.53 ;
        RECT 2.4 -4.16 2.5 -3.625 ;
        RECT 2.4 -2.835 2.5 -2.3 ;
        RECT 2.4 -0.93 2.5 -0.395 ;
        RECT 2.4 0.395 2.5 0.93 ;
        RECT 1.2 -49.38 1.3 -48.845 ;
        RECT 1.2 -48.055 1.3 -47.52 ;
        RECT 1.2 -46.15 1.3 -45.615 ;
        RECT 1.2 -44.825 1.3 -44.29 ;
        RECT 1.2 -42.92 1.3 -42.385 ;
        RECT 1.2 -41.595 1.3 -41.06 ;
        RECT 1.2 -39.69 1.3 -39.155 ;
        RECT 1.2 -38.365 1.3 -37.83 ;
        RECT 1.2 -36.46 1.3 -35.925 ;
        RECT 1.2 -35.135 1.3 -34.6 ;
        RECT 1.2 -33.23 1.3 -32.695 ;
        RECT 1.2 -31.905 1.3 -31.37 ;
        RECT 1.2 -30 1.3 -29.465 ;
        RECT 1.2 -28.675 1.3 -28.14 ;
        RECT 1.2 -26.77 1.3 -26.235 ;
        RECT 1.2 -25.445 1.3 -24.91 ;
        RECT 1.2 -23.54 1.3 -23.005 ;
        RECT 1.2 -22.215 1.3 -21.68 ;
        RECT 1.2 -20.31 1.3 -19.775 ;
        RECT 1.2 -18.985 1.3 -18.45 ;
        RECT 1.2 -17.08 1.3 -16.545 ;
        RECT 1.2 -15.755 1.3 -15.22 ;
        RECT 1.2 -13.85 1.3 -13.315 ;
        RECT 1.2 -12.525 1.3 -11.99 ;
        RECT 1.2 -10.62 1.3 -10.085 ;
        RECT 1.2 -9.295 1.3 -8.76 ;
        RECT 1.2 -7.39 1.3 -6.855 ;
        RECT 1.2 -6.065 1.3 -5.53 ;
        RECT 1.2 -4.16 1.3 -3.625 ;
        RECT 1.2 -2.835 1.3 -2.3 ;
        RECT 1.2 -0.93 1.3 -0.395 ;
        RECT 1.2 0.395 1.3 0.93 ;
        RECT 0 -49.38 0.1 -48.845 ;
        RECT 0 -48.055 0.1 -47.52 ;
        RECT 0 -46.15 0.1 -45.615 ;
        RECT 0 -44.825 0.1 -44.29 ;
        RECT 0 -42.92 0.1 -42.385 ;
        RECT 0 -41.595 0.1 -41.06 ;
        RECT 0 -39.69 0.1 -39.155 ;
        RECT 0 -38.365 0.1 -37.83 ;
        RECT 0 -36.46 0.1 -35.925 ;
        RECT 0 -35.135 0.1 -34.6 ;
        RECT 0 -33.23 0.1 -32.695 ;
        RECT 0 -31.905 0.1 -31.37 ;
        RECT 0 -30 0.1 -29.465 ;
        RECT 0 -28.675 0.1 -28.14 ;
        RECT 0 -26.77 0.1 -26.235 ;
        RECT 0 -25.445 0.1 -24.91 ;
        RECT 0 -23.54 0.1 -23.005 ;
        RECT 0 -22.215 0.1 -21.68 ;
        RECT 0 -20.31 0.1 -19.775 ;
        RECT 0 -18.985 0.1 -18.45 ;
        RECT 0 -17.08 0.1 -16.545 ;
        RECT 0 -15.755 0.1 -15.22 ;
        RECT 0 -13.85 0.1 -13.315 ;
        RECT 0 -12.525 0.1 -11.99 ;
        RECT 0 -10.62 0.1 -10.085 ;
        RECT 0 -9.295 0.1 -8.76 ;
        RECT 0 -7.39 0.1 -6.855 ;
        RECT 0 -6.065 0.1 -5.53 ;
        RECT 0 -4.16 0.1 -3.625 ;
        RECT 0 -2.835 0.1 -2.3 ;
        RECT 0 -0.93 0.1 -0.395 ;
        RECT 0 0.395 0.1 0.93 ;
        RECT -33.525 -56.865 -0.585 -56.185 ;
        RECT -1.025 -56.865 -0.925 -55.555 ;
        RECT -1.805 -56.865 -1.705 -55.375 ;
        RECT -2.325 -56.865 -2.225 -55.555 ;
        RECT -3.105 -56.865 -3.005 -55.375 ;
        RECT -3.625 -56.865 -3.525 -55.555 ;
        RECT -4.405 -56.865 -4.305 -55.375 ;
        RECT -4.925 -56.865 -4.825 -55.555 ;
        RECT -5.705 -56.865 -5.605 -55.375 ;
        RECT -6.225 -56.865 -6.125 -55.555 ;
        RECT -7.005 -56.865 -6.905 -55.375 ;
        RECT -7.525 -56.865 -7.425 -55.555 ;
        RECT -8.305 -56.865 -8.205 -55.375 ;
        RECT -8.825 -56.865 -8.725 -55.555 ;
        RECT -9.605 -56.865 -9.505 -55.375 ;
        RECT -10.125 -56.865 -10.025 -55.555 ;
        RECT -10.905 -56.865 -10.805 -55.375 ;
        RECT -11.525 -57.495 -11.425 -56.185 ;
        RECT -12.125 -57.495 -12.025 -56.185 ;
        RECT -33.525 -43.945 -0.585 -43.265 ;
        RECT -1.025 -44.575 -0.925 -42.635 ;
        RECT -1.805 -44.755 -1.705 -42.455 ;
        RECT -2.325 -44.575 -2.225 -42.635 ;
        RECT -3.105 -44.755 -3.005 -42.455 ;
        RECT -3.625 -44.575 -3.525 -42.635 ;
        RECT -4.405 -44.755 -4.305 -42.455 ;
        RECT -4.925 -44.575 -4.825 -42.635 ;
        RECT -5.705 -44.755 -5.605 -42.455 ;
        RECT -6.225 -44.575 -6.125 -42.635 ;
        RECT -7.005 -44.755 -6.905 -42.455 ;
        RECT -7.525 -44.575 -7.425 -42.635 ;
        RECT -8.305 -44.755 -8.205 -42.455 ;
        RECT -8.825 -44.575 -8.725 -42.635 ;
        RECT -9.605 -44.755 -9.505 -42.455 ;
        RECT -10.125 -44.575 -10.025 -42.635 ;
        RECT -10.905 -44.755 -10.805 -42.455 ;
        RECT -11.425 -44.575 -11.325 -42.635 ;
        RECT -12.205 -44.755 -12.105 -42.455 ;
        RECT -12.725 -44.575 -12.625 -42.635 ;
        RECT -13.505 -44.755 -13.405 -42.455 ;
        RECT -14.025 -44.575 -13.925 -42.635 ;
        RECT -14.805 -44.755 -14.705 -42.455 ;
        RECT -15.325 -44.575 -15.225 -42.635 ;
        RECT -16.105 -44.755 -16.005 -42.455 ;
        RECT -16.625 -44.575 -16.525 -42.635 ;
        RECT -17.405 -44.755 -17.305 -42.455 ;
        RECT -17.925 -44.575 -17.825 -42.635 ;
        RECT -18.705 -44.755 -18.605 -42.455 ;
        RECT -19.225 -44.575 -19.125 -42.635 ;
        RECT -20.005 -44.755 -19.905 -42.455 ;
        RECT -20.525 -44.575 -20.425 -42.635 ;
        RECT -21.305 -44.755 -21.205 -42.455 ;
        RECT -21.825 -44.575 -21.725 -42.635 ;
        RECT -22.605 -44.755 -22.505 -42.455 ;
        RECT -23.125 -44.575 -23.025 -42.635 ;
        RECT -23.905 -44.755 -23.805 -42.455 ;
        RECT -24.425 -44.575 -24.325 -42.635 ;
        RECT -25.205 -44.755 -25.105 -42.455 ;
        RECT -25.725 -44.575 -25.625 -42.635 ;
        RECT -26.505 -44.755 -26.405 -42.455 ;
        RECT -33.525 -31.025 -0.585 -30.345 ;
        RECT -1.025 -31.655 -0.925 -29.715 ;
        RECT -1.805 -31.835 -1.705 -29.535 ;
        RECT -2.325 -31.655 -2.225 -29.715 ;
        RECT -3.105 -31.835 -3.005 -29.535 ;
        RECT -3.625 -31.655 -3.525 -29.715 ;
        RECT -4.405 -31.835 -4.305 -29.535 ;
        RECT -4.925 -31.655 -4.825 -29.715 ;
        RECT -5.705 -31.835 -5.605 -29.535 ;
        RECT -6.225 -31.655 -6.125 -29.715 ;
        RECT -7.005 -31.835 -6.905 -29.535 ;
        RECT -7.525 -31.655 -7.425 -29.715 ;
        RECT -8.305 -31.835 -8.205 -29.535 ;
        RECT -8.825 -31.655 -8.725 -29.715 ;
        RECT -9.605 -31.835 -9.505 -29.535 ;
        RECT -10.125 -31.655 -10.025 -29.715 ;
        RECT -10.905 -31.835 -10.805 -29.535 ;
        RECT -11.425 -31.655 -11.325 -29.715 ;
        RECT -12.205 -31.835 -12.105 -29.535 ;
        RECT -12.725 -31.655 -12.625 -29.715 ;
        RECT -13.505 -31.835 -13.405 -29.535 ;
        RECT -14.025 -31.655 -13.925 -29.715 ;
        RECT -14.805 -31.835 -14.705 -29.535 ;
        RECT -15.325 -31.655 -15.225 -29.715 ;
        RECT -16.105 -31.835 -16.005 -29.535 ;
        RECT -16.625 -31.655 -16.525 -29.715 ;
        RECT -17.405 -31.835 -17.305 -29.535 ;
        RECT -17.925 -31.655 -17.825 -29.715 ;
        RECT -18.705 -31.835 -18.605 -29.535 ;
        RECT -19.225 -31.655 -19.125 -29.715 ;
        RECT -20.005 -31.835 -19.905 -29.535 ;
        RECT -20.525 -31.655 -20.425 -29.715 ;
        RECT -21.305 -31.835 -21.205 -29.535 ;
        RECT -21.825 -31.655 -21.725 -29.715 ;
        RECT -22.605 -31.835 -22.505 -29.535 ;
        RECT -23.125 -31.655 -23.025 -29.715 ;
        RECT -23.905 -31.835 -23.805 -29.535 ;
        RECT -24.425 -31.655 -24.325 -29.715 ;
        RECT -25.205 -31.835 -25.105 -29.535 ;
        RECT -25.725 -31.655 -25.625 -29.715 ;
        RECT -26.505 -31.835 -26.405 -29.535 ;
        RECT -33.525 -18.105 -0.585 -17.425 ;
        RECT -1.025 -18.735 -0.925 -16.795 ;
        RECT -1.805 -18.915 -1.705 -16.615 ;
        RECT -2.325 -18.735 -2.225 -16.795 ;
        RECT -3.105 -18.915 -3.005 -16.615 ;
        RECT -3.625 -18.735 -3.525 -16.795 ;
        RECT -4.405 -18.915 -4.305 -16.615 ;
        RECT -4.925 -18.735 -4.825 -16.795 ;
        RECT -5.705 -18.915 -5.605 -16.615 ;
        RECT -6.225 -18.735 -6.125 -16.795 ;
        RECT -7.005 -18.915 -6.905 -16.615 ;
        RECT -7.525 -18.735 -7.425 -16.795 ;
        RECT -8.305 -18.915 -8.205 -16.615 ;
        RECT -8.825 -18.735 -8.725 -16.795 ;
        RECT -9.605 -18.915 -9.505 -16.615 ;
        RECT -10.125 -18.735 -10.025 -16.795 ;
        RECT -10.905 -18.915 -10.805 -16.615 ;
        RECT -11.425 -18.735 -11.325 -16.795 ;
        RECT -12.205 -18.915 -12.105 -16.615 ;
        RECT -12.725 -18.735 -12.625 -16.795 ;
        RECT -13.505 -18.915 -13.405 -16.615 ;
        RECT -14.025 -18.735 -13.925 -16.795 ;
        RECT -14.805 -18.915 -14.705 -16.615 ;
        RECT -15.325 -18.735 -15.225 -16.795 ;
        RECT -16.105 -18.915 -16.005 -16.615 ;
        RECT -16.625 -18.735 -16.525 -16.795 ;
        RECT -17.405 -18.915 -17.305 -16.615 ;
        RECT -17.925 -18.735 -17.825 -16.795 ;
        RECT -18.705 -18.915 -18.605 -16.615 ;
        RECT -19.225 -18.735 -19.125 -16.795 ;
        RECT -20.005 -18.915 -19.905 -16.615 ;
        RECT -20.525 -18.735 -20.425 -16.795 ;
        RECT -21.305 -18.915 -21.205 -16.615 ;
        RECT -21.825 -18.735 -21.725 -16.795 ;
        RECT -22.605 -18.915 -22.505 -16.615 ;
        RECT -23.125 -18.735 -23.025 -16.795 ;
        RECT -23.905 -18.915 -23.805 -16.615 ;
        RECT -24.425 -18.735 -24.325 -16.795 ;
        RECT -25.205 -18.915 -25.105 -16.615 ;
        RECT -25.725 -18.735 -25.625 -16.795 ;
        RECT -26.505 -18.915 -26.405 -16.615 ;
        RECT -33.525 -5.185 -0.585 -4.505 ;
        RECT -1.025 -5.815 -0.925 -3.875 ;
        RECT -1.805 -5.995 -1.705 -3.695 ;
        RECT -2.325 -5.815 -2.225 -3.875 ;
        RECT -3.105 -5.995 -3.005 -3.695 ;
        RECT -3.625 -5.815 -3.525 -3.875 ;
        RECT -4.405 -5.995 -4.305 -3.695 ;
        RECT -4.925 -5.815 -4.825 -3.875 ;
        RECT -5.705 -5.995 -5.605 -3.695 ;
        RECT -6.225 -5.815 -6.125 -3.875 ;
        RECT -7.005 -5.995 -6.905 -3.695 ;
        RECT -7.525 -5.815 -7.425 -3.875 ;
        RECT -8.305 -5.995 -8.205 -3.695 ;
        RECT -8.825 -5.815 -8.725 -3.875 ;
        RECT -9.605 -5.995 -9.505 -3.695 ;
        RECT -10.125 -5.815 -10.025 -3.875 ;
        RECT -10.905 -5.995 -10.805 -3.695 ;
        RECT -11.425 -5.815 -11.325 -3.875 ;
        RECT -12.205 -5.995 -12.105 -3.695 ;
        RECT -12.725 -5.815 -12.625 -3.875 ;
        RECT -13.505 -5.995 -13.405 -3.695 ;
        RECT -14.025 -5.815 -13.925 -3.875 ;
        RECT -14.805 -5.995 -14.705 -3.695 ;
        RECT -15.325 -5.815 -15.225 -3.875 ;
        RECT -16.105 -5.995 -16.005 -3.695 ;
        RECT -16.625 -5.815 -16.525 -3.875 ;
        RECT -17.405 -5.995 -17.305 -3.695 ;
        RECT -17.925 -5.815 -17.825 -3.875 ;
        RECT -18.705 -5.995 -18.605 -3.695 ;
        RECT -19.225 -5.815 -19.125 -3.875 ;
        RECT -20.005 -5.995 -19.905 -3.695 ;
        RECT -20.525 -5.815 -20.425 -3.875 ;
        RECT -21.305 -5.995 -21.205 -3.695 ;
        RECT -21.825 -5.815 -21.725 -3.875 ;
        RECT -22.605 -5.995 -22.505 -3.695 ;
        RECT -23.125 -5.815 -23.025 -3.875 ;
        RECT -23.905 -5.995 -23.805 -3.695 ;
        RECT -24.425 -5.815 -24.325 -3.875 ;
        RECT -25.205 -5.995 -25.105 -3.695 ;
        RECT -25.725 -5.815 -25.625 -3.875 ;
        RECT -26.505 -5.995 -26.405 -3.695 ;
        RECT -33.525 5.275 -26.565 5.955 ;
        RECT -27.125 4.645 -27.025 5.955 ;
        RECT -27.725 4.645 -27.625 5.955 ;
        RECT -28.325 4.645 -28.225 5.955 ;
        RECT -28.925 4.645 -28.825 5.955 ;
        RECT -29.525 4.645 -29.425 5.955 ;
        RECT 0.025 -63.775 43.265 -63.415 ;
        RECT 34.64 -63.775 34.74 -63 ;
        RECT 34.08 -63.775 34.18 -63 ;
        RECT 29.84 -63.775 29.94 -63 ;
        RECT 29.28 -63.775 29.38 -63 ;
        RECT 25.04 -63.775 25.14 -63 ;
        RECT 24.48 -63.775 24.58 -63 ;
        RECT 20.24 -63.775 20.34 -63 ;
        RECT 19.68 -63.775 19.78 -63 ;
        RECT 15.44 -63.775 15.54 -63 ;
        RECT 14.88 -63.775 14.98 -63 ;
        RECT 10.64 -63.775 10.74 -63 ;
        RECT 10.08 -63.775 10.18 -63 ;
        RECT 5.84 -63.775 5.94 -63 ;
        RECT 5.28 -63.775 5.38 -63 ;
        RECT 1.04 -63.775 1.14 -63 ;
        RECT 0.48 -63.775 0.58 -63 ;
        RECT 0.01 -58.515 43.265 -58.155 ;
        RECT 38.005 -59.085 38.105 -58.155 ;
        RECT 37.675 -58.515 37.775 -57.59 ;
        RECT 37.445 -59.085 37.545 -58.155 ;
        RECT 37.115 -58.515 37.215 -57.59 ;
        RECT 36.295 -59.07 36.395 -58.155 ;
        RECT 35.985 -59.085 36.085 -58.155 ;
        RECT 35.675 -58.515 35.775 -57.59 ;
        RECT 35.425 -59.085 35.525 -58.155 ;
        RECT 35.115 -58.515 35.215 -57.59 ;
        RECT 34.24 -59.085 34.415 -58.155 ;
        RECT 33.685 -59.05 33.785 -58.155 ;
        RECT 33.205 -59.085 33.305 -58.155 ;
        RECT 32.875 -58.515 32.975 -57.59 ;
        RECT 32.645 -59.085 32.745 -58.155 ;
        RECT 32.315 -58.515 32.415 -57.59 ;
        RECT 31.495 -59.07 31.595 -58.155 ;
        RECT 31.185 -59.085 31.285 -58.155 ;
        RECT 30.875 -58.515 30.975 -57.59 ;
        RECT 30.625 -59.085 30.725 -58.155 ;
        RECT 30.315 -58.515 30.415 -57.59 ;
        RECT 29.44 -59.085 29.615 -58.155 ;
        RECT 28.885 -59.05 28.985 -58.155 ;
        RECT 28.405 -59.085 28.505 -58.155 ;
        RECT 28.075 -58.515 28.175 -57.59 ;
        RECT 27.845 -59.085 27.945 -58.155 ;
        RECT 27.515 -58.515 27.615 -57.59 ;
        RECT 26.695 -59.07 26.795 -58.155 ;
        RECT 26.385 -59.085 26.485 -58.155 ;
        RECT 26.075 -58.515 26.175 -57.59 ;
        RECT 25.825 -59.085 25.925 -58.155 ;
        RECT 25.515 -58.515 25.615 -57.59 ;
        RECT 24.64 -59.085 24.815 -58.155 ;
        RECT 24.085 -59.05 24.185 -58.155 ;
        RECT 23.605 -59.085 23.705 -58.155 ;
        RECT 23.275 -58.515 23.375 -57.59 ;
        RECT 23.045 -59.085 23.145 -58.155 ;
        RECT 22.715 -58.515 22.815 -57.59 ;
        RECT 21.895 -59.07 21.995 -58.155 ;
        RECT 21.585 -59.085 21.685 -58.155 ;
        RECT 21.275 -58.515 21.375 -57.59 ;
        RECT 21.025 -59.085 21.125 -58.155 ;
        RECT 20.715 -58.515 20.815 -57.59 ;
        RECT 19.84 -59.085 20.015 -58.155 ;
        RECT 19.285 -59.05 19.385 -58.155 ;
        RECT 18.805 -59.085 18.905 -58.155 ;
        RECT 18.475 -58.515 18.575 -57.59 ;
        RECT 18.245 -59.085 18.345 -58.155 ;
        RECT 17.915 -58.515 18.015 -57.59 ;
        RECT 17.095 -59.07 17.195 -58.155 ;
        RECT 16.785 -59.085 16.885 -58.155 ;
        RECT 16.475 -58.515 16.575 -57.59 ;
        RECT 16.225 -59.085 16.325 -58.155 ;
        RECT 15.915 -58.515 16.015 -57.59 ;
        RECT 15.04 -59.085 15.215 -58.155 ;
        RECT 14.485 -59.05 14.585 -58.155 ;
        RECT 14.005 -59.085 14.105 -58.155 ;
        RECT 13.675 -58.515 13.775 -57.59 ;
        RECT 13.445 -59.085 13.545 -58.155 ;
        RECT 13.115 -58.515 13.215 -57.59 ;
        RECT 12.295 -59.07 12.395 -58.155 ;
        RECT 11.985 -59.085 12.085 -58.155 ;
        RECT 11.675 -58.515 11.775 -57.59 ;
        RECT 11.425 -59.085 11.525 -58.155 ;
        RECT 11.115 -58.515 11.215 -57.59 ;
        RECT 10.24 -59.085 10.415 -58.155 ;
        RECT 9.685 -59.05 9.785 -58.155 ;
        RECT 9.205 -59.085 9.305 -58.155 ;
        RECT 8.875 -58.515 8.975 -57.59 ;
        RECT 8.645 -59.085 8.745 -58.155 ;
        RECT 8.315 -58.515 8.415 -57.59 ;
        RECT 7.495 -59.07 7.595 -58.155 ;
        RECT 7.185 -59.085 7.285 -58.155 ;
        RECT 6.875 -58.515 6.975 -57.59 ;
        RECT 6.625 -59.085 6.725 -58.155 ;
        RECT 6.315 -58.515 6.415 -57.59 ;
        RECT 5.44 -59.085 5.615 -58.155 ;
        RECT 4.885 -59.05 4.985 -58.155 ;
        RECT 4.405 -59.085 4.505 -58.155 ;
        RECT 4.075 -58.515 4.175 -57.59 ;
        RECT 3.845 -59.085 3.945 -58.155 ;
        RECT 3.515 -58.515 3.615 -57.59 ;
        RECT 2.695 -59.07 2.795 -58.155 ;
        RECT 2.385 -59.085 2.485 -58.155 ;
        RECT 2.075 -58.515 2.175 -57.59 ;
        RECT 1.825 -59.085 1.925 -58.155 ;
        RECT 1.515 -58.515 1.615 -57.59 ;
        RECT 0.64 -59.085 0.815 -58.155 ;
        RECT 0.085 -59.05 0.185 -58.155 ;
        RECT -33.525 7.175 43.265 9.895 ;
        RECT -6.48 4.965 -5.245 9.895 ;
        RECT -5.885 4.385 -5.785 9.895 ;
        RECT 38.4 -49.38 38.5 -48.845 ;
        RECT 38.4 -48.055 38.5 -47.52 ;
        RECT 38.4 -46.15 38.5 -45.615 ;
        RECT 38.4 -44.825 38.5 -44.29 ;
        RECT 38.4 -42.92 38.5 -42.385 ;
        RECT 38.4 -41.595 38.5 -41.06 ;
        RECT 38.4 -39.69 38.5 -39.155 ;
        RECT 38.4 -38.365 38.5 -37.83 ;
        RECT 38.4 -36.46 38.5 -35.925 ;
        RECT 38.4 -35.135 38.5 -34.6 ;
        RECT 38.4 -33.23 38.5 -32.695 ;
        RECT 38.4 -31.905 38.5 -31.37 ;
        RECT 38.4 -30 38.5 -29.465 ;
        RECT 38.4 -28.675 38.5 -28.14 ;
        RECT 38.4 -26.77 38.5 -26.235 ;
        RECT 38.4 -25.445 38.5 -24.91 ;
        RECT 38.4 -23.54 38.5 -23.005 ;
        RECT 38.4 -22.215 38.5 -21.68 ;
        RECT 38.4 -20.31 38.5 -19.775 ;
        RECT 38.4 -18.985 38.5 -18.45 ;
        RECT 38.4 -17.08 38.5 -16.545 ;
        RECT 38.4 -15.755 38.5 -15.22 ;
        RECT 38.4 -13.85 38.5 -13.315 ;
        RECT 38.4 -12.525 38.5 -11.99 ;
        RECT 38.4 -10.62 38.5 -10.085 ;
        RECT 38.4 -9.295 38.5 -8.76 ;
        RECT 38.4 -7.39 38.5 -6.855 ;
        RECT 38.4 -6.065 38.5 -5.53 ;
        RECT 38.4 -4.16 38.5 -3.625 ;
        RECT 38.4 -2.835 38.5 -2.3 ;
        RECT 38.4 -0.93 38.5 -0.395 ;
        RECT 38.4 0.395 38.5 0.93 ;
        RECT 37.2 -49.38 37.3 -48.845 ;
        RECT 37.2 -48.055 37.3 -47.52 ;
        RECT 37.2 -46.15 37.3 -45.615 ;
        RECT 37.2 -44.825 37.3 -44.29 ;
        RECT 37.2 -42.92 37.3 -42.385 ;
        RECT 37.2 -41.595 37.3 -41.06 ;
        RECT 37.2 -39.69 37.3 -39.155 ;
        RECT 37.2 -38.365 37.3 -37.83 ;
        RECT 37.2 -36.46 37.3 -35.925 ;
        RECT 37.2 -35.135 37.3 -34.6 ;
        RECT 37.2 -33.23 37.3 -32.695 ;
        RECT 37.2 -31.905 37.3 -31.37 ;
        RECT 37.2 -30 37.3 -29.465 ;
        RECT 37.2 -28.675 37.3 -28.14 ;
        RECT 37.2 -26.77 37.3 -26.235 ;
        RECT 37.2 -25.445 37.3 -24.91 ;
        RECT 37.2 -23.54 37.3 -23.005 ;
        RECT 37.2 -22.215 37.3 -21.68 ;
        RECT 37.2 -20.31 37.3 -19.775 ;
        RECT 37.2 -18.985 37.3 -18.45 ;
        RECT 37.2 -17.08 37.3 -16.545 ;
        RECT 37.2 -15.755 37.3 -15.22 ;
        RECT 37.2 -13.85 37.3 -13.315 ;
        RECT 37.2 -12.525 37.3 -11.99 ;
        RECT 37.2 -10.62 37.3 -10.085 ;
        RECT 37.2 -9.295 37.3 -8.76 ;
        RECT 37.2 -7.39 37.3 -6.855 ;
        RECT 37.2 -6.065 37.3 -5.53 ;
        RECT 37.2 -4.16 37.3 -3.625 ;
        RECT 37.2 -2.835 37.3 -2.3 ;
        RECT 37.2 -0.93 37.3 -0.395 ;
        RECT 37.2 0.395 37.3 0.93 ;
        RECT 36 -49.38 36.1 -48.845 ;
        RECT 36 -48.055 36.1 -47.52 ;
        RECT 36 -46.15 36.1 -45.615 ;
        RECT 36 -44.825 36.1 -44.29 ;
        RECT 36 -42.92 36.1 -42.385 ;
        RECT 36 -41.595 36.1 -41.06 ;
        RECT 36 -39.69 36.1 -39.155 ;
        RECT 36 -38.365 36.1 -37.83 ;
        RECT 36 -36.46 36.1 -35.925 ;
        RECT 36 -35.135 36.1 -34.6 ;
        RECT 36 -33.23 36.1 -32.695 ;
        RECT 36 -31.905 36.1 -31.37 ;
        RECT 36 -30 36.1 -29.465 ;
        RECT 36 -28.675 36.1 -28.14 ;
        RECT 36 -26.77 36.1 -26.235 ;
        RECT 36 -25.445 36.1 -24.91 ;
        RECT 36 -23.54 36.1 -23.005 ;
        RECT 36 -22.215 36.1 -21.68 ;
        RECT 36 -20.31 36.1 -19.775 ;
        RECT 36 -18.985 36.1 -18.45 ;
        RECT 36 -17.08 36.1 -16.545 ;
        RECT 36 -15.755 36.1 -15.22 ;
        RECT 36 -13.85 36.1 -13.315 ;
        RECT 36 -12.525 36.1 -11.99 ;
        RECT 36 -10.62 36.1 -10.085 ;
        RECT 36 -9.295 36.1 -8.76 ;
        RECT 36 -7.39 36.1 -6.855 ;
        RECT 36 -6.065 36.1 -5.53 ;
        RECT 36 -4.16 36.1 -3.625 ;
        RECT 36 -2.835 36.1 -2.3 ;
        RECT 36 -0.93 36.1 -0.395 ;
        RECT 36 0.395 36.1 0.93 ;
        RECT 34.8 -49.38 34.9 -48.845 ;
        RECT 34.8 -48.055 34.9 -47.52 ;
        RECT 34.8 -46.15 34.9 -45.615 ;
        RECT 34.8 -44.825 34.9 -44.29 ;
        RECT 34.8 -42.92 34.9 -42.385 ;
        RECT 34.8 -41.595 34.9 -41.06 ;
        RECT 34.8 -39.69 34.9 -39.155 ;
        RECT 34.8 -38.365 34.9 -37.83 ;
        RECT 34.8 -36.46 34.9 -35.925 ;
        RECT 34.8 -35.135 34.9 -34.6 ;
        RECT 34.8 -33.23 34.9 -32.695 ;
        RECT 34.8 -31.905 34.9 -31.37 ;
        RECT 34.8 -30 34.9 -29.465 ;
        RECT 34.8 -28.675 34.9 -28.14 ;
        RECT 34.8 -26.77 34.9 -26.235 ;
        RECT 34.8 -25.445 34.9 -24.91 ;
        RECT 34.8 -23.54 34.9 -23.005 ;
        RECT 34.8 -22.215 34.9 -21.68 ;
        RECT 34.8 -20.31 34.9 -19.775 ;
        RECT 34.8 -18.985 34.9 -18.45 ;
        RECT 34.8 -17.08 34.9 -16.545 ;
        RECT 34.8 -15.755 34.9 -15.22 ;
        RECT 34.8 -13.85 34.9 -13.315 ;
        RECT 34.8 -12.525 34.9 -11.99 ;
        RECT 34.8 -10.62 34.9 -10.085 ;
        RECT 34.8 -9.295 34.9 -8.76 ;
        RECT 34.8 -7.39 34.9 -6.855 ;
        RECT 34.8 -6.065 34.9 -5.53 ;
        RECT 34.8 -4.16 34.9 -3.625 ;
        RECT 34.8 -2.835 34.9 -2.3 ;
        RECT 34.8 -0.93 34.9 -0.395 ;
        RECT 34.8 0.395 34.9 0.93 ;
        RECT 33.6 -49.38 33.7 -48.845 ;
        RECT 33.6 -48.055 33.7 -47.52 ;
        RECT 33.6 -46.15 33.7 -45.615 ;
        RECT 33.6 -44.825 33.7 -44.29 ;
        RECT 33.6 -42.92 33.7 -42.385 ;
        RECT 33.6 -41.595 33.7 -41.06 ;
        RECT 33.6 -39.69 33.7 -39.155 ;
        RECT 33.6 -38.365 33.7 -37.83 ;
        RECT 33.6 -36.46 33.7 -35.925 ;
        RECT 33.6 -35.135 33.7 -34.6 ;
        RECT 33.6 -33.23 33.7 -32.695 ;
        RECT 33.6 -31.905 33.7 -31.37 ;
        RECT 33.6 -30 33.7 -29.465 ;
        RECT 33.6 -28.675 33.7 -28.14 ;
        RECT 33.6 -26.77 33.7 -26.235 ;
        RECT 33.6 -25.445 33.7 -24.91 ;
        RECT 33.6 -23.54 33.7 -23.005 ;
        RECT 33.6 -22.215 33.7 -21.68 ;
        RECT 33.6 -20.31 33.7 -19.775 ;
        RECT 33.6 -18.985 33.7 -18.45 ;
        RECT 33.6 -17.08 33.7 -16.545 ;
        RECT 33.6 -15.755 33.7 -15.22 ;
        RECT 33.6 -13.85 33.7 -13.315 ;
        RECT 33.6 -12.525 33.7 -11.99 ;
        RECT 33.6 -10.62 33.7 -10.085 ;
        RECT 33.6 -9.295 33.7 -8.76 ;
        RECT 33.6 -7.39 33.7 -6.855 ;
        RECT 33.6 -6.065 33.7 -5.53 ;
        RECT 33.6 -4.16 33.7 -3.625 ;
        RECT 33.6 -2.835 33.7 -2.3 ;
        RECT 33.6 -0.93 33.7 -0.395 ;
        RECT 33.6 0.395 33.7 0.93 ;
        RECT 32.4 -49.38 32.5 -48.845 ;
        RECT 32.4 -48.055 32.5 -47.52 ;
        RECT 32.4 -46.15 32.5 -45.615 ;
        RECT 32.4 -44.825 32.5 -44.29 ;
        RECT 32.4 -42.92 32.5 -42.385 ;
        RECT 32.4 -41.595 32.5 -41.06 ;
        RECT 32.4 -39.69 32.5 -39.155 ;
        RECT 32.4 -38.365 32.5 -37.83 ;
        RECT 32.4 -36.46 32.5 -35.925 ;
        RECT 32.4 -35.135 32.5 -34.6 ;
        RECT 32.4 -33.23 32.5 -32.695 ;
        RECT 32.4 -31.905 32.5 -31.37 ;
        RECT 32.4 -30 32.5 -29.465 ;
        RECT 32.4 -28.675 32.5 -28.14 ;
        RECT 32.4 -26.77 32.5 -26.235 ;
        RECT 32.4 -25.445 32.5 -24.91 ;
        RECT 32.4 -23.54 32.5 -23.005 ;
        RECT 32.4 -22.215 32.5 -21.68 ;
        RECT 32.4 -20.31 32.5 -19.775 ;
        RECT 32.4 -18.985 32.5 -18.45 ;
        RECT 32.4 -17.08 32.5 -16.545 ;
        RECT 32.4 -15.755 32.5 -15.22 ;
        RECT 32.4 -13.85 32.5 -13.315 ;
        RECT 32.4 -12.525 32.5 -11.99 ;
        RECT 32.4 -10.62 32.5 -10.085 ;
        RECT 32.4 -9.295 32.5 -8.76 ;
        RECT 32.4 -7.39 32.5 -6.855 ;
        RECT 32.4 -6.065 32.5 -5.53 ;
        RECT 32.4 -4.16 32.5 -3.625 ;
        RECT 32.4 -2.835 32.5 -2.3 ;
        RECT 32.4 -0.93 32.5 -0.395 ;
        RECT 32.4 0.395 32.5 0.93 ;
        RECT 31.2 -49.38 31.3 -48.845 ;
        RECT 31.2 -48.055 31.3 -47.52 ;
        RECT 31.2 -46.15 31.3 -45.615 ;
        RECT 31.2 -44.825 31.3 -44.29 ;
        RECT 31.2 -42.92 31.3 -42.385 ;
        RECT 31.2 -41.595 31.3 -41.06 ;
        RECT 31.2 -39.69 31.3 -39.155 ;
        RECT 31.2 -38.365 31.3 -37.83 ;
        RECT 31.2 -36.46 31.3 -35.925 ;
        RECT 31.2 -35.135 31.3 -34.6 ;
        RECT 31.2 -33.23 31.3 -32.695 ;
        RECT 31.2 -31.905 31.3 -31.37 ;
        RECT 31.2 -30 31.3 -29.465 ;
        RECT 31.2 -28.675 31.3 -28.14 ;
        RECT 31.2 -26.77 31.3 -26.235 ;
        RECT 31.2 -25.445 31.3 -24.91 ;
        RECT 31.2 -23.54 31.3 -23.005 ;
        RECT 31.2 -22.215 31.3 -21.68 ;
        RECT 31.2 -20.31 31.3 -19.775 ;
        RECT 31.2 -18.985 31.3 -18.45 ;
        RECT 31.2 -17.08 31.3 -16.545 ;
        RECT 31.2 -15.755 31.3 -15.22 ;
        RECT 31.2 -13.85 31.3 -13.315 ;
        RECT 31.2 -12.525 31.3 -11.99 ;
        RECT 31.2 -10.62 31.3 -10.085 ;
        RECT 31.2 -9.295 31.3 -8.76 ;
        RECT 31.2 -7.39 31.3 -6.855 ;
        RECT 31.2 -6.065 31.3 -5.53 ;
        RECT 31.2 -4.16 31.3 -3.625 ;
        RECT 31.2 -2.835 31.3 -2.3 ;
        RECT 31.2 -0.93 31.3 -0.395 ;
        RECT 31.2 0.395 31.3 0.93 ;
        RECT 30 -49.38 30.1 -48.845 ;
        RECT 30 -48.055 30.1 -47.52 ;
        RECT 30 -46.15 30.1 -45.615 ;
        RECT 30 -44.825 30.1 -44.29 ;
        RECT 30 -42.92 30.1 -42.385 ;
        RECT 30 -41.595 30.1 -41.06 ;
        RECT 30 -39.69 30.1 -39.155 ;
        RECT 30 -38.365 30.1 -37.83 ;
        RECT 30 -36.46 30.1 -35.925 ;
        RECT 30 -35.135 30.1 -34.6 ;
        RECT 30 -33.23 30.1 -32.695 ;
        RECT 30 -31.905 30.1 -31.37 ;
        RECT 30 -30 30.1 -29.465 ;
        RECT 30 -28.675 30.1 -28.14 ;
        RECT 30 -26.77 30.1 -26.235 ;
        RECT 30 -25.445 30.1 -24.91 ;
        RECT 30 -23.54 30.1 -23.005 ;
        RECT 30 -22.215 30.1 -21.68 ;
        RECT 30 -20.31 30.1 -19.775 ;
        RECT 30 -18.985 30.1 -18.45 ;
        RECT 30 -17.08 30.1 -16.545 ;
        RECT 30 -15.755 30.1 -15.22 ;
        RECT 30 -13.85 30.1 -13.315 ;
        RECT 30 -12.525 30.1 -11.99 ;
        RECT 30 -10.62 30.1 -10.085 ;
        RECT 30 -9.295 30.1 -8.76 ;
        RECT 30 -7.39 30.1 -6.855 ;
        RECT 30 -6.065 30.1 -5.53 ;
        RECT 30 -4.16 30.1 -3.625 ;
        RECT 30 -2.835 30.1 -2.3 ;
        RECT 30 -0.93 30.1 -0.395 ;
        RECT 30 0.395 30.1 0.93 ;
        RECT 28.8 -49.38 28.9 -48.845 ;
        RECT 28.8 -48.055 28.9 -47.52 ;
        RECT 28.8 -46.15 28.9 -45.615 ;
        RECT 28.8 -44.825 28.9 -44.29 ;
        RECT 28.8 -42.92 28.9 -42.385 ;
        RECT 28.8 -41.595 28.9 -41.06 ;
        RECT 28.8 -39.69 28.9 -39.155 ;
        RECT 28.8 -38.365 28.9 -37.83 ;
        RECT 28.8 -36.46 28.9 -35.925 ;
        RECT 28.8 -35.135 28.9 -34.6 ;
        RECT 28.8 -33.23 28.9 -32.695 ;
        RECT 28.8 -31.905 28.9 -31.37 ;
        RECT 28.8 -30 28.9 -29.465 ;
        RECT 28.8 -28.675 28.9 -28.14 ;
        RECT 28.8 -26.77 28.9 -26.235 ;
        RECT 28.8 -25.445 28.9 -24.91 ;
        RECT 28.8 -23.54 28.9 -23.005 ;
        RECT 28.8 -22.215 28.9 -21.68 ;
        RECT 28.8 -20.31 28.9 -19.775 ;
        RECT 28.8 -18.985 28.9 -18.45 ;
        RECT 28.8 -17.08 28.9 -16.545 ;
        RECT 28.8 -15.755 28.9 -15.22 ;
        RECT 28.8 -13.85 28.9 -13.315 ;
        RECT 28.8 -12.525 28.9 -11.99 ;
        RECT 28.8 -10.62 28.9 -10.085 ;
        RECT 28.8 -9.295 28.9 -8.76 ;
        RECT 28.8 -7.39 28.9 -6.855 ;
        RECT 28.8 -6.065 28.9 -5.53 ;
        RECT 28.8 -4.16 28.9 -3.625 ;
        RECT 28.8 -2.835 28.9 -2.3 ;
        RECT 28.8 -0.93 28.9 -0.395 ;
        RECT 28.8 0.395 28.9 0.93 ;
        RECT 27.6 -49.38 27.7 -48.845 ;
        RECT 27.6 -48.055 27.7 -47.52 ;
        RECT 27.6 -46.15 27.7 -45.615 ;
        RECT 27.6 -44.825 27.7 -44.29 ;
        RECT 27.6 -42.92 27.7 -42.385 ;
        RECT 27.6 -41.595 27.7 -41.06 ;
        RECT 27.6 -39.69 27.7 -39.155 ;
        RECT 27.6 -38.365 27.7 -37.83 ;
        RECT 27.6 -36.46 27.7 -35.925 ;
        RECT 27.6 -35.135 27.7 -34.6 ;
        RECT 27.6 -33.23 27.7 -32.695 ;
        RECT 27.6 -31.905 27.7 -31.37 ;
        RECT 27.6 -30 27.7 -29.465 ;
        RECT 27.6 -28.675 27.7 -28.14 ;
        RECT 27.6 -26.77 27.7 -26.235 ;
        RECT 27.6 -25.445 27.7 -24.91 ;
        RECT 27.6 -23.54 27.7 -23.005 ;
        RECT 27.6 -22.215 27.7 -21.68 ;
        RECT 27.6 -20.31 27.7 -19.775 ;
        RECT 27.6 -18.985 27.7 -18.45 ;
        RECT 27.6 -17.08 27.7 -16.545 ;
        RECT 27.6 -15.755 27.7 -15.22 ;
        RECT 27.6 -13.85 27.7 -13.315 ;
        RECT 27.6 -12.525 27.7 -11.99 ;
        RECT 27.6 -10.62 27.7 -10.085 ;
        RECT 27.6 -9.295 27.7 -8.76 ;
        RECT 27.6 -7.39 27.7 -6.855 ;
        RECT 27.6 -6.065 27.7 -5.53 ;
        RECT 27.6 -4.16 27.7 -3.625 ;
        RECT 27.6 -2.835 27.7 -2.3 ;
        RECT 27.6 -0.93 27.7 -0.395 ;
        RECT 27.6 0.395 27.7 0.93 ;
        RECT 26.4 -49.38 26.5 -48.845 ;
        RECT 26.4 -48.055 26.5 -47.52 ;
        RECT 26.4 -46.15 26.5 -45.615 ;
        RECT 26.4 -44.825 26.5 -44.29 ;
        RECT 26.4 -42.92 26.5 -42.385 ;
        RECT 26.4 -41.595 26.5 -41.06 ;
        RECT 26.4 -39.69 26.5 -39.155 ;
        RECT 26.4 -38.365 26.5 -37.83 ;
        RECT 26.4 -36.46 26.5 -35.925 ;
        RECT 26.4 -35.135 26.5 -34.6 ;
        RECT 26.4 -33.23 26.5 -32.695 ;
        RECT 26.4 -31.905 26.5 -31.37 ;
        RECT 26.4 -30 26.5 -29.465 ;
        RECT 26.4 -28.675 26.5 -28.14 ;
        RECT 26.4 -26.77 26.5 -26.235 ;
        RECT 26.4 -25.445 26.5 -24.91 ;
        RECT 26.4 -23.54 26.5 -23.005 ;
        RECT 26.4 -22.215 26.5 -21.68 ;
        RECT 26.4 -20.31 26.5 -19.775 ;
        RECT 26.4 -18.985 26.5 -18.45 ;
        RECT 26.4 -17.08 26.5 -16.545 ;
        RECT 26.4 -15.755 26.5 -15.22 ;
        RECT 26.4 -13.85 26.5 -13.315 ;
        RECT 26.4 -12.525 26.5 -11.99 ;
        RECT 26.4 -10.62 26.5 -10.085 ;
        RECT 26.4 -9.295 26.5 -8.76 ;
        RECT 26.4 -7.39 26.5 -6.855 ;
        RECT 26.4 -6.065 26.5 -5.53 ;
        RECT 26.4 -4.16 26.5 -3.625 ;
        RECT 26.4 -2.835 26.5 -2.3 ;
        RECT 26.4 -0.93 26.5 -0.395 ;
        RECT 26.4 0.395 26.5 0.93 ;
        RECT 25.2 -49.38 25.3 -48.845 ;
        RECT 25.2 -48.055 25.3 -47.52 ;
        RECT 25.2 -46.15 25.3 -45.615 ;
        RECT 25.2 -44.825 25.3 -44.29 ;
        RECT 25.2 -42.92 25.3 -42.385 ;
        RECT 25.2 -41.595 25.3 -41.06 ;
        RECT 25.2 -39.69 25.3 -39.155 ;
        RECT 25.2 -38.365 25.3 -37.83 ;
        RECT 25.2 -36.46 25.3 -35.925 ;
        RECT 25.2 -35.135 25.3 -34.6 ;
        RECT 25.2 -33.23 25.3 -32.695 ;
        RECT 25.2 -31.905 25.3 -31.37 ;
        RECT 25.2 -30 25.3 -29.465 ;
        RECT 25.2 -28.675 25.3 -28.14 ;
        RECT 25.2 -26.77 25.3 -26.235 ;
        RECT 25.2 -25.445 25.3 -24.91 ;
        RECT 25.2 -23.54 25.3 -23.005 ;
        RECT 25.2 -22.215 25.3 -21.68 ;
        RECT 25.2 -20.31 25.3 -19.775 ;
        RECT 25.2 -18.985 25.3 -18.45 ;
        RECT 25.2 -17.08 25.3 -16.545 ;
        RECT 25.2 -15.755 25.3 -15.22 ;
        RECT 25.2 -13.85 25.3 -13.315 ;
        RECT 25.2 -12.525 25.3 -11.99 ;
        RECT 25.2 -10.62 25.3 -10.085 ;
        RECT 25.2 -9.295 25.3 -8.76 ;
        RECT 25.2 -7.39 25.3 -6.855 ;
        RECT 25.2 -6.065 25.3 -5.53 ;
        RECT 25.2 -4.16 25.3 -3.625 ;
        RECT 25.2 -2.835 25.3 -2.3 ;
        RECT 25.2 -0.93 25.3 -0.395 ;
        RECT 25.2 0.395 25.3 0.93 ;
        RECT 24 -49.38 24.1 -48.845 ;
        RECT 24 -48.055 24.1 -47.52 ;
        RECT 24 -46.15 24.1 -45.615 ;
        RECT 24 -44.825 24.1 -44.29 ;
        RECT 24 -42.92 24.1 -42.385 ;
        RECT 24 -41.595 24.1 -41.06 ;
        RECT 24 -39.69 24.1 -39.155 ;
        RECT 24 -38.365 24.1 -37.83 ;
        RECT 24 -36.46 24.1 -35.925 ;
        RECT 24 -35.135 24.1 -34.6 ;
        RECT 24 -33.23 24.1 -32.695 ;
        RECT 24 -31.905 24.1 -31.37 ;
        RECT 24 -30 24.1 -29.465 ;
        RECT 24 -28.675 24.1 -28.14 ;
        RECT 24 -26.77 24.1 -26.235 ;
        RECT 24 -25.445 24.1 -24.91 ;
        RECT 24 -23.54 24.1 -23.005 ;
        RECT 24 -22.215 24.1 -21.68 ;
        RECT 24 -20.31 24.1 -19.775 ;
        RECT 24 -18.985 24.1 -18.45 ;
        RECT 24 -17.08 24.1 -16.545 ;
        RECT 24 -15.755 24.1 -15.22 ;
        RECT 24 -13.85 24.1 -13.315 ;
        RECT 24 -12.525 24.1 -11.99 ;
        RECT 24 -10.62 24.1 -10.085 ;
        RECT 24 -9.295 24.1 -8.76 ;
        RECT 24 -7.39 24.1 -6.855 ;
        RECT 24 -6.065 24.1 -5.53 ;
        RECT 24 -4.16 24.1 -3.625 ;
        RECT 24 -2.835 24.1 -2.3 ;
        RECT 24 -0.93 24.1 -0.395 ;
        RECT 24 0.395 24.1 0.93 ;
        RECT 22.8 -49.38 22.9 -48.845 ;
        RECT 22.8 -48.055 22.9 -47.52 ;
        RECT 22.8 -46.15 22.9 -45.615 ;
        RECT 22.8 -44.825 22.9 -44.29 ;
        RECT 22.8 -42.92 22.9 -42.385 ;
        RECT 22.8 -41.595 22.9 -41.06 ;
        RECT 22.8 -39.69 22.9 -39.155 ;
        RECT 22.8 -38.365 22.9 -37.83 ;
        RECT 22.8 -36.46 22.9 -35.925 ;
        RECT 22.8 -35.135 22.9 -34.6 ;
        RECT 22.8 -33.23 22.9 -32.695 ;
        RECT 22.8 -31.905 22.9 -31.37 ;
        RECT 22.8 -30 22.9 -29.465 ;
        RECT 22.8 -28.675 22.9 -28.14 ;
        RECT 22.8 -26.77 22.9 -26.235 ;
        RECT 22.8 -25.445 22.9 -24.91 ;
        RECT 22.8 -23.54 22.9 -23.005 ;
        RECT 22.8 -22.215 22.9 -21.68 ;
        RECT 22.8 -20.31 22.9 -19.775 ;
        RECT 22.8 -18.985 22.9 -18.45 ;
        RECT 22.8 -17.08 22.9 -16.545 ;
        RECT 22.8 -15.755 22.9 -15.22 ;
        RECT 22.8 -13.85 22.9 -13.315 ;
        RECT 22.8 -12.525 22.9 -11.99 ;
        RECT 22.8 -10.62 22.9 -10.085 ;
        RECT 22.8 -9.295 22.9 -8.76 ;
        RECT 22.8 -7.39 22.9 -6.855 ;
        RECT 22.8 -6.065 22.9 -5.53 ;
        RECT 22.8 -4.16 22.9 -3.625 ;
        RECT 22.8 -2.835 22.9 -2.3 ;
        RECT 22.8 -0.93 22.9 -0.395 ;
        RECT 22.8 0.395 22.9 0.93 ;
        RECT 21.6 -49.38 21.7 -48.845 ;
        RECT 21.6 -48.055 21.7 -47.52 ;
        RECT 21.6 -46.15 21.7 -45.615 ;
        RECT 21.6 -44.825 21.7 -44.29 ;
        RECT 21.6 -42.92 21.7 -42.385 ;
        RECT 21.6 -41.595 21.7 -41.06 ;
        RECT 21.6 -39.69 21.7 -39.155 ;
        RECT 21.6 -38.365 21.7 -37.83 ;
        RECT 21.6 -36.46 21.7 -35.925 ;
        RECT 21.6 -35.135 21.7 -34.6 ;
        RECT 21.6 -33.23 21.7 -32.695 ;
        RECT 21.6 -31.905 21.7 -31.37 ;
        RECT 21.6 -30 21.7 -29.465 ;
        RECT 21.6 -28.675 21.7 -28.14 ;
        RECT 21.6 -26.77 21.7 -26.235 ;
        RECT 21.6 -25.445 21.7 -24.91 ;
        RECT 21.6 -23.54 21.7 -23.005 ;
        RECT 21.6 -22.215 21.7 -21.68 ;
        RECT 21.6 -20.31 21.7 -19.775 ;
        RECT 21.6 -18.985 21.7 -18.45 ;
        RECT 21.6 -17.08 21.7 -16.545 ;
        RECT 21.6 -15.755 21.7 -15.22 ;
        RECT 21.6 -13.85 21.7 -13.315 ;
        RECT 21.6 -12.525 21.7 -11.99 ;
        RECT 21.6 -10.62 21.7 -10.085 ;
        RECT 21.6 -9.295 21.7 -8.76 ;
        RECT 21.6 -7.39 21.7 -6.855 ;
        RECT 21.6 -6.065 21.7 -5.53 ;
        RECT 21.6 -4.16 21.7 -3.625 ;
        RECT 21.6 -2.835 21.7 -2.3 ;
        RECT 21.6 -0.93 21.7 -0.395 ;
        RECT 21.6 0.395 21.7 0.93 ;
        RECT 20.4 -49.38 20.5 -48.845 ;
        RECT 20.4 -48.055 20.5 -47.52 ;
        RECT 20.4 -46.15 20.5 -45.615 ;
        RECT 20.4 -44.825 20.5 -44.29 ;
        RECT 20.4 -42.92 20.5 -42.385 ;
        RECT 20.4 -41.595 20.5 -41.06 ;
        RECT 20.4 -39.69 20.5 -39.155 ;
        RECT 20.4 -38.365 20.5 -37.83 ;
        RECT 20.4 -36.46 20.5 -35.925 ;
        RECT 20.4 -35.135 20.5 -34.6 ;
        RECT 20.4 -33.23 20.5 -32.695 ;
        RECT 20.4 -31.905 20.5 -31.37 ;
        RECT 20.4 -30 20.5 -29.465 ;
        RECT 20.4 -28.675 20.5 -28.14 ;
        RECT 20.4 -26.77 20.5 -26.235 ;
        RECT 20.4 -25.445 20.5 -24.91 ;
        RECT 20.4 -23.54 20.5 -23.005 ;
        RECT 20.4 -22.215 20.5 -21.68 ;
        RECT 20.4 -20.31 20.5 -19.775 ;
        RECT 20.4 -18.985 20.5 -18.45 ;
        RECT 20.4 -17.08 20.5 -16.545 ;
        RECT 20.4 -15.755 20.5 -15.22 ;
        RECT 20.4 -13.85 20.5 -13.315 ;
        RECT 20.4 -12.525 20.5 -11.99 ;
        RECT 20.4 -10.62 20.5 -10.085 ;
        RECT 20.4 -9.295 20.5 -8.76 ;
        RECT 20.4 -7.39 20.5 -6.855 ;
        RECT 20.4 -6.065 20.5 -5.53 ;
        RECT 20.4 -4.16 20.5 -3.625 ;
        RECT 20.4 -2.835 20.5 -2.3 ;
        RECT 20.4 -0.93 20.5 -0.395 ;
        RECT 20.4 0.395 20.5 0.93 ;
        RECT 19.2 -49.38 19.3 -48.845 ;
        RECT 19.2 -48.055 19.3 -47.52 ;
        RECT 19.2 -46.15 19.3 -45.615 ;
        RECT 19.2 -44.825 19.3 -44.29 ;
        RECT 19.2 -42.92 19.3 -42.385 ;
        RECT 19.2 -41.595 19.3 -41.06 ;
        RECT 19.2 -39.69 19.3 -39.155 ;
        RECT 19.2 -38.365 19.3 -37.83 ;
        RECT 19.2 -36.46 19.3 -35.925 ;
        RECT 19.2 -35.135 19.3 -34.6 ;
        RECT 19.2 -33.23 19.3 -32.695 ;
        RECT 19.2 -31.905 19.3 -31.37 ;
        RECT 19.2 -30 19.3 -29.465 ;
        RECT 19.2 -28.675 19.3 -28.14 ;
        RECT 19.2 -26.77 19.3 -26.235 ;
        RECT 19.2 -25.445 19.3 -24.91 ;
        RECT 19.2 -23.54 19.3 -23.005 ;
        RECT 19.2 -22.215 19.3 -21.68 ;
        RECT 19.2 -20.31 19.3 -19.775 ;
        RECT 19.2 -18.985 19.3 -18.45 ;
        RECT 19.2 -17.08 19.3 -16.545 ;
        RECT 19.2 -15.755 19.3 -15.22 ;
        RECT 19.2 -13.85 19.3 -13.315 ;
        RECT 19.2 -12.525 19.3 -11.99 ;
        RECT 19.2 -10.62 19.3 -10.085 ;
        RECT 19.2 -9.295 19.3 -8.76 ;
        RECT 19.2 -7.39 19.3 -6.855 ;
        RECT 19.2 -6.065 19.3 -5.53 ;
        RECT 19.2 -4.16 19.3 -3.625 ;
        RECT 19.2 -2.835 19.3 -2.3 ;
        RECT 19.2 -0.93 19.3 -0.395 ;
        RECT 19.2 0.395 19.3 0.93 ;
        RECT 18 -49.38 18.1 -48.845 ;
        RECT 18 -48.055 18.1 -47.52 ;
        RECT 18 -46.15 18.1 -45.615 ;
        RECT 18 -44.825 18.1 -44.29 ;
        RECT 18 -42.92 18.1 -42.385 ;
        RECT 18 -41.595 18.1 -41.06 ;
        RECT 18 -39.69 18.1 -39.155 ;
        RECT 18 -38.365 18.1 -37.83 ;
        RECT 18 -36.46 18.1 -35.925 ;
        RECT 18 -35.135 18.1 -34.6 ;
        RECT 18 -33.23 18.1 -32.695 ;
        RECT 18 -31.905 18.1 -31.37 ;
        RECT 18 -30 18.1 -29.465 ;
        RECT 18 -28.675 18.1 -28.14 ;
        RECT 18 -26.77 18.1 -26.235 ;
        RECT 18 -25.445 18.1 -24.91 ;
        RECT 18 -23.54 18.1 -23.005 ;
        RECT 18 -22.215 18.1 -21.68 ;
        RECT 18 -20.31 18.1 -19.775 ;
        RECT 18 -18.985 18.1 -18.45 ;
        RECT 18 -17.08 18.1 -16.545 ;
        RECT 18 -15.755 18.1 -15.22 ;
        RECT 18 -13.85 18.1 -13.315 ;
        RECT 18 -12.525 18.1 -11.99 ;
        RECT 18 -10.62 18.1 -10.085 ;
        RECT 18 -9.295 18.1 -8.76 ;
        RECT 18 -7.39 18.1 -6.855 ;
        RECT 18 -6.065 18.1 -5.53 ;
        RECT 18 -4.16 18.1 -3.625 ;
        RECT 18 -2.835 18.1 -2.3 ;
        RECT 18 -0.93 18.1 -0.395 ;
        RECT 18 0.395 18.1 0.93 ;
        RECT 16.8 -49.38 16.9 -48.845 ;
        RECT 16.8 -48.055 16.9 -47.52 ;
        RECT 16.8 -46.15 16.9 -45.615 ;
        RECT 16.8 -44.825 16.9 -44.29 ;
        RECT 16.8 -42.92 16.9 -42.385 ;
        RECT 16.8 -41.595 16.9 -41.06 ;
        RECT 16.8 -39.69 16.9 -39.155 ;
        RECT 16.8 -38.365 16.9 -37.83 ;
        RECT 16.8 -36.46 16.9 -35.925 ;
        RECT 16.8 -35.135 16.9 -34.6 ;
        RECT 16.8 -33.23 16.9 -32.695 ;
        RECT 16.8 -31.905 16.9 -31.37 ;
        RECT 16.8 -30 16.9 -29.465 ;
        RECT 16.8 -28.675 16.9 -28.14 ;
        RECT 16.8 -26.77 16.9 -26.235 ;
        RECT 16.8 -25.445 16.9 -24.91 ;
        RECT 16.8 -23.54 16.9 -23.005 ;
        RECT 16.8 -22.215 16.9 -21.68 ;
        RECT 16.8 -20.31 16.9 -19.775 ;
        RECT 16.8 -18.985 16.9 -18.45 ;
        RECT 16.8 -17.08 16.9 -16.545 ;
        RECT 16.8 -15.755 16.9 -15.22 ;
        RECT 16.8 -13.85 16.9 -13.315 ;
        RECT 16.8 -12.525 16.9 -11.99 ;
        RECT 16.8 -10.62 16.9 -10.085 ;
        RECT 16.8 -9.295 16.9 -8.76 ;
        RECT 16.8 -7.39 16.9 -6.855 ;
        RECT 16.8 -6.065 16.9 -5.53 ;
        RECT 16.8 -4.16 16.9 -3.625 ;
        RECT 16.8 -2.835 16.9 -2.3 ;
        RECT 16.8 -0.93 16.9 -0.395 ;
        RECT 16.8 0.395 16.9 0.93 ;
        RECT 15.6 -49.38 15.7 -48.845 ;
        RECT 15.6 -48.055 15.7 -47.52 ;
        RECT 15.6 -46.15 15.7 -45.615 ;
        RECT 15.6 -44.825 15.7 -44.29 ;
        RECT 15.6 -42.92 15.7 -42.385 ;
        RECT 15.6 -41.595 15.7 -41.06 ;
        RECT 15.6 -39.69 15.7 -39.155 ;
        RECT 15.6 -38.365 15.7 -37.83 ;
        RECT 15.6 -36.46 15.7 -35.925 ;
        RECT 15.6 -35.135 15.7 -34.6 ;
        RECT 15.6 -33.23 15.7 -32.695 ;
        RECT 15.6 -31.905 15.7 -31.37 ;
        RECT 15.6 -30 15.7 -29.465 ;
        RECT 15.6 -28.675 15.7 -28.14 ;
        RECT 15.6 -26.77 15.7 -26.235 ;
        RECT 15.6 -25.445 15.7 -24.91 ;
        RECT 15.6 -23.54 15.7 -23.005 ;
        RECT 15.6 -22.215 15.7 -21.68 ;
        RECT 15.6 -20.31 15.7 -19.775 ;
        RECT 15.6 -18.985 15.7 -18.45 ;
        RECT 15.6 -17.08 15.7 -16.545 ;
        RECT 15.6 -15.755 15.7 -15.22 ;
        RECT 15.6 -13.85 15.7 -13.315 ;
        RECT 15.6 -12.525 15.7 -11.99 ;
        RECT 15.6 -10.62 15.7 -10.085 ;
        RECT 15.6 -9.295 15.7 -8.76 ;
        RECT 15.6 -7.39 15.7 -6.855 ;
        RECT 15.6 -6.065 15.7 -5.53 ;
        RECT 15.6 -4.16 15.7 -3.625 ;
        RECT 15.6 -2.835 15.7 -2.3 ;
        RECT 15.6 -0.93 15.7 -0.395 ;
        RECT 15.6 0.395 15.7 0.93 ;
        RECT 14.4 -49.38 14.5 -48.845 ;
        RECT 14.4 -48.055 14.5 -47.52 ;
        RECT 14.4 -46.15 14.5 -45.615 ;
        RECT 14.4 -44.825 14.5 -44.29 ;
        RECT 14.4 -42.92 14.5 -42.385 ;
        RECT 14.4 -41.595 14.5 -41.06 ;
        RECT 14.4 -39.69 14.5 -39.155 ;
        RECT 14.4 -38.365 14.5 -37.83 ;
        RECT 14.4 -36.46 14.5 -35.925 ;
        RECT 14.4 -35.135 14.5 -34.6 ;
        RECT 14.4 -33.23 14.5 -32.695 ;
        RECT 14.4 -31.905 14.5 -31.37 ;
        RECT 14.4 -30 14.5 -29.465 ;
        RECT 14.4 -28.675 14.5 -28.14 ;
        RECT 14.4 -26.77 14.5 -26.235 ;
        RECT 14.4 -25.445 14.5 -24.91 ;
        RECT 14.4 -23.54 14.5 -23.005 ;
        RECT 14.4 -22.215 14.5 -21.68 ;
        RECT 14.4 -20.31 14.5 -19.775 ;
        RECT 14.4 -18.985 14.5 -18.45 ;
        RECT 14.4 -17.08 14.5 -16.545 ;
        RECT 14.4 -15.755 14.5 -15.22 ;
        RECT 14.4 -13.85 14.5 -13.315 ;
        RECT 14.4 -12.525 14.5 -11.99 ;
        RECT 14.4 -10.62 14.5 -10.085 ;
        RECT 14.4 -9.295 14.5 -8.76 ;
        RECT 14.4 -7.39 14.5 -6.855 ;
        RECT 14.4 -6.065 14.5 -5.53 ;
        RECT 14.4 -4.16 14.5 -3.625 ;
        RECT 14.4 -2.835 14.5 -2.3 ;
        RECT 14.4 -0.93 14.5 -0.395 ;
        RECT 14.4 0.395 14.5 0.93 ;
        RECT 13.2 -49.38 13.3 -48.845 ;
        RECT 13.2 -48.055 13.3 -47.52 ;
        RECT 13.2 -46.15 13.3 -45.615 ;
        RECT 13.2 -44.825 13.3 -44.29 ;
        RECT 13.2 -42.92 13.3 -42.385 ;
        RECT 13.2 -41.595 13.3 -41.06 ;
        RECT 13.2 -39.69 13.3 -39.155 ;
        RECT 13.2 -38.365 13.3 -37.83 ;
        RECT 13.2 -36.46 13.3 -35.925 ;
        RECT 13.2 -35.135 13.3 -34.6 ;
        RECT 13.2 -33.23 13.3 -32.695 ;
        RECT 13.2 -31.905 13.3 -31.37 ;
        RECT 13.2 -30 13.3 -29.465 ;
        RECT 13.2 -28.675 13.3 -28.14 ;
        RECT 13.2 -26.77 13.3 -26.235 ;
        RECT 13.2 -25.445 13.3 -24.91 ;
        RECT 13.2 -23.54 13.3 -23.005 ;
        RECT 13.2 -22.215 13.3 -21.68 ;
        RECT 13.2 -20.31 13.3 -19.775 ;
        RECT 13.2 -18.985 13.3 -18.45 ;
        RECT 13.2 -17.08 13.3 -16.545 ;
        RECT 13.2 -15.755 13.3 -15.22 ;
        RECT 13.2 -13.85 13.3 -13.315 ;
        RECT 13.2 -12.525 13.3 -11.99 ;
        RECT 13.2 -10.62 13.3 -10.085 ;
        RECT 13.2 -9.295 13.3 -8.76 ;
        RECT 13.2 -7.39 13.3 -6.855 ;
        RECT 13.2 -6.065 13.3 -5.53 ;
        RECT 13.2 -4.16 13.3 -3.625 ;
        RECT 13.2 -2.835 13.3 -2.3 ;
        RECT 13.2 -0.93 13.3 -0.395 ;
        RECT 13.2 0.395 13.3 0.93 ;
        RECT 12 -49.38 12.1 -48.845 ;
        RECT 12 -48.055 12.1 -47.52 ;
        RECT 12 -46.15 12.1 -45.615 ;
        RECT 12 -44.825 12.1 -44.29 ;
        RECT 12 -42.92 12.1 -42.385 ;
        RECT 12 -41.595 12.1 -41.06 ;
        RECT 12 -39.69 12.1 -39.155 ;
        RECT 12 -38.365 12.1 -37.83 ;
        RECT 12 -36.46 12.1 -35.925 ;
        RECT 12 -35.135 12.1 -34.6 ;
        RECT 12 -33.23 12.1 -32.695 ;
        RECT 12 -31.905 12.1 -31.37 ;
        RECT 12 -30 12.1 -29.465 ;
        RECT 12 -28.675 12.1 -28.14 ;
        RECT 12 -26.77 12.1 -26.235 ;
        RECT 12 -25.445 12.1 -24.91 ;
        RECT 12 -23.54 12.1 -23.005 ;
        RECT 12 -22.215 12.1 -21.68 ;
        RECT 12 -20.31 12.1 -19.775 ;
        RECT 12 -18.985 12.1 -18.45 ;
        RECT 12 -17.08 12.1 -16.545 ;
        RECT 12 -15.755 12.1 -15.22 ;
        RECT 12 -13.85 12.1 -13.315 ;
        RECT 12 -12.525 12.1 -11.99 ;
        RECT 12 -10.62 12.1 -10.085 ;
        RECT 12 -9.295 12.1 -8.76 ;
        RECT 12 -7.39 12.1 -6.855 ;
        RECT 12 -6.065 12.1 -5.53 ;
        RECT 12 -4.16 12.1 -3.625 ;
        RECT 12 -2.835 12.1 -2.3 ;
        RECT 12 -0.93 12.1 -0.395 ;
        RECT 12 0.395 12.1 0.93 ;
        RECT 10.8 -49.38 10.9 -48.845 ;
        RECT 10.8 -48.055 10.9 -47.52 ;
        RECT 10.8 -46.15 10.9 -45.615 ;
        RECT 10.8 -44.825 10.9 -44.29 ;
        RECT 10.8 -42.92 10.9 -42.385 ;
        RECT 10.8 -41.595 10.9 -41.06 ;
        RECT 10.8 -39.69 10.9 -39.155 ;
        RECT 10.8 -38.365 10.9 -37.83 ;
        RECT 10.8 -36.46 10.9 -35.925 ;
        RECT 10.8 -35.135 10.9 -34.6 ;
        RECT 10.8 -33.23 10.9 -32.695 ;
        RECT 10.8 -31.905 10.9 -31.37 ;
        RECT 10.8 -30 10.9 -29.465 ;
        RECT 10.8 -28.675 10.9 -28.14 ;
        RECT 10.8 -26.77 10.9 -26.235 ;
        RECT 10.8 -25.445 10.9 -24.91 ;
        RECT 10.8 -23.54 10.9 -23.005 ;
        RECT 10.8 -22.215 10.9 -21.68 ;
        RECT 10.8 -20.31 10.9 -19.775 ;
        RECT 10.8 -18.985 10.9 -18.45 ;
        RECT 10.8 -17.08 10.9 -16.545 ;
        RECT 10.8 -15.755 10.9 -15.22 ;
        RECT 10.8 -13.85 10.9 -13.315 ;
        RECT 10.8 -12.525 10.9 -11.99 ;
        RECT 10.8 -10.62 10.9 -10.085 ;
        RECT 10.8 -9.295 10.9 -8.76 ;
        RECT 10.8 -7.39 10.9 -6.855 ;
        RECT 10.8 -6.065 10.9 -5.53 ;
        RECT 10.8 -4.16 10.9 -3.625 ;
        RECT 10.8 -2.835 10.9 -2.3 ;
        RECT 10.8 -0.93 10.9 -0.395 ;
        RECT 10.8 0.395 10.9 0.93 ;
        RECT 9.6 -49.38 9.7 -48.845 ;
        RECT 9.6 -48.055 9.7 -47.52 ;
        RECT 9.6 -46.15 9.7 -45.615 ;
        RECT 9.6 -44.825 9.7 -44.29 ;
        RECT 9.6 -42.92 9.7 -42.385 ;
        RECT 9.6 -41.595 9.7 -41.06 ;
        RECT 9.6 -39.69 9.7 -39.155 ;
        RECT 9.6 -38.365 9.7 -37.83 ;
        RECT 9.6 -36.46 9.7 -35.925 ;
        RECT 9.6 -35.135 9.7 -34.6 ;
        RECT 9.6 -33.23 9.7 -32.695 ;
        RECT 9.6 -31.905 9.7 -31.37 ;
        RECT 9.6 -30 9.7 -29.465 ;
        RECT 9.6 -28.675 9.7 -28.14 ;
        RECT 9.6 -26.77 9.7 -26.235 ;
        RECT 9.6 -25.445 9.7 -24.91 ;
        RECT 9.6 -23.54 9.7 -23.005 ;
        RECT 9.6 -22.215 9.7 -21.68 ;
        RECT 9.6 -20.31 9.7 -19.775 ;
        RECT 9.6 -18.985 9.7 -18.45 ;
        RECT 9.6 -17.08 9.7 -16.545 ;
        RECT 9.6 -15.755 9.7 -15.22 ;
        RECT 9.6 -13.85 9.7 -13.315 ;
        RECT 9.6 -12.525 9.7 -11.99 ;
        RECT 9.6 -10.62 9.7 -10.085 ;
        RECT 9.6 -9.295 9.7 -8.76 ;
        RECT 9.6 -7.39 9.7 -6.855 ;
        RECT 9.6 -6.065 9.7 -5.53 ;
        RECT 9.6 -4.16 9.7 -3.625 ;
        RECT 9.6 -2.835 9.7 -2.3 ;
        RECT 9.6 -0.93 9.7 -0.395 ;
        RECT 9.6 0.395 9.7 0.93 ;
        RECT 8.4 -49.38 8.5 -48.845 ;
        RECT 8.4 -48.055 8.5 -47.52 ;
        RECT 8.4 -46.15 8.5 -45.615 ;
        RECT 8.4 -44.825 8.5 -44.29 ;
        RECT 8.4 -42.92 8.5 -42.385 ;
        RECT 8.4 -41.595 8.5 -41.06 ;
        RECT 8.4 -39.69 8.5 -39.155 ;
        RECT 8.4 -38.365 8.5 -37.83 ;
        RECT 8.4 -36.46 8.5 -35.925 ;
        RECT 8.4 -35.135 8.5 -34.6 ;
        RECT 8.4 -33.23 8.5 -32.695 ;
        RECT 8.4 -31.905 8.5 -31.37 ;
        RECT 8.4 -30 8.5 -29.465 ;
        RECT 8.4 -28.675 8.5 -28.14 ;
        RECT 8.4 -26.77 8.5 -26.235 ;
        RECT 8.4 -25.445 8.5 -24.91 ;
        RECT 8.4 -23.54 8.5 -23.005 ;
        RECT 8.4 -22.215 8.5 -21.68 ;
        RECT 8.4 -20.31 8.5 -19.775 ;
        RECT 8.4 -18.985 8.5 -18.45 ;
        RECT 8.4 -17.08 8.5 -16.545 ;
        RECT 8.4 -15.755 8.5 -15.22 ;
        RECT 8.4 -13.85 8.5 -13.315 ;
        RECT 8.4 -12.525 8.5 -11.99 ;
        RECT 8.4 -10.62 8.5 -10.085 ;
        RECT 8.4 -9.295 8.5 -8.76 ;
        RECT 8.4 -7.39 8.5 -6.855 ;
        RECT 8.4 -6.065 8.5 -5.53 ;
        RECT 8.4 -4.16 8.5 -3.625 ;
        RECT 8.4 -2.835 8.5 -2.3 ;
        RECT 8.4 -0.93 8.5 -0.395 ;
        RECT 8.4 0.395 8.5 0.93 ;
        RECT 7.2 -49.38 7.3 -48.845 ;
        RECT 7.2 -48.055 7.3 -47.52 ;
        RECT 7.2 -46.15 7.3 -45.615 ;
        RECT 7.2 -44.825 7.3 -44.29 ;
        RECT 7.2 -42.92 7.3 -42.385 ;
        RECT 7.2 -41.595 7.3 -41.06 ;
        RECT 7.2 -39.69 7.3 -39.155 ;
        RECT 7.2 -38.365 7.3 -37.83 ;
        RECT 7.2 -36.46 7.3 -35.925 ;
        RECT 7.2 -35.135 7.3 -34.6 ;
        RECT 7.2 -33.23 7.3 -32.695 ;
        RECT 7.2 -31.905 7.3 -31.37 ;
        RECT 7.2 -30 7.3 -29.465 ;
        RECT 7.2 -28.675 7.3 -28.14 ;
        RECT 7.2 -26.77 7.3 -26.235 ;
        RECT 7.2 -25.445 7.3 -24.91 ;
        RECT 7.2 -23.54 7.3 -23.005 ;
        RECT 7.2 -22.215 7.3 -21.68 ;
        RECT 7.2 -20.31 7.3 -19.775 ;
        RECT 7.2 -18.985 7.3 -18.45 ;
        RECT 7.2 -17.08 7.3 -16.545 ;
        RECT 7.2 -15.755 7.3 -15.22 ;
        RECT 7.2 -13.85 7.3 -13.315 ;
        RECT 7.2 -12.525 7.3 -11.99 ;
        RECT 7.2 -10.62 7.3 -10.085 ;
        RECT 7.2 -9.295 7.3 -8.76 ;
        RECT 7.2 -7.39 7.3 -6.855 ;
        RECT 7.2 -6.065 7.3 -5.53 ;
        RECT 7.2 -4.16 7.3 -3.625 ;
        RECT 7.2 -2.835 7.3 -2.3 ;
        RECT 7.2 -0.93 7.3 -0.395 ;
        RECT 7.2 0.395 7.3 0.93 ;
        RECT 6 -49.38 6.1 -48.845 ;
        RECT 6 -48.055 6.1 -47.52 ;
        RECT 6 -46.15 6.1 -45.615 ;
        RECT 6 -44.825 6.1 -44.29 ;
        RECT 6 -42.92 6.1 -42.385 ;
        RECT 6 -41.595 6.1 -41.06 ;
        RECT 6 -39.69 6.1 -39.155 ;
        RECT 6 -38.365 6.1 -37.83 ;
        RECT 6 -36.46 6.1 -35.925 ;
        RECT 6 -35.135 6.1 -34.6 ;
        RECT 6 -33.23 6.1 -32.695 ;
        RECT 6 -31.905 6.1 -31.37 ;
        RECT 6 -30 6.1 -29.465 ;
        RECT 6 -28.675 6.1 -28.14 ;
        RECT 6 -26.77 6.1 -26.235 ;
        RECT 6 -25.445 6.1 -24.91 ;
        RECT 6 -23.54 6.1 -23.005 ;
        RECT 6 -22.215 6.1 -21.68 ;
        RECT 6 -20.31 6.1 -19.775 ;
        RECT 6 -18.985 6.1 -18.45 ;
        RECT 6 -17.08 6.1 -16.545 ;
        RECT 6 -15.755 6.1 -15.22 ;
        RECT 6 -13.85 6.1 -13.315 ;
        RECT 6 -12.525 6.1 -11.99 ;
        RECT 6 -10.62 6.1 -10.085 ;
        RECT 6 -9.295 6.1 -8.76 ;
        RECT 6 -7.39 6.1 -6.855 ;
      LAYER V1 ;
        RECT 27.6 -37.96 27.7 -37.86 ;
        RECT 27.6 -38.315 27.7 -38.215 ;
        RECT 27.6 -39.305 27.7 -39.205 ;
        RECT 27.6 -39.66 27.7 -39.56 ;
        RECT 27.6 -41.19 27.7 -41.09 ;
        RECT 27.6 -41.545 27.7 -41.445 ;
        RECT 27.6 -42.535 27.7 -42.435 ;
        RECT 27.6 -42.89 27.7 -42.79 ;
        RECT 27.6 -44.42 27.7 -44.32 ;
        RECT 27.6 -44.775 27.7 -44.675 ;
        RECT 27.6 -45.765 27.7 -45.665 ;
        RECT 27.6 -46.12 27.7 -46.02 ;
        RECT 27.6 -47.65 27.7 -47.55 ;
        RECT 27.6 -48.005 27.7 -47.905 ;
        RECT 27.6 -48.995 27.7 -48.895 ;
        RECT 27.6 -49.35 27.7 -49.25 ;
        RECT 28.8 9.75 28.9 9.85 ;
        RECT 28.8 9.52 28.9 9.62 ;
        RECT 28.8 9.29 28.9 9.39 ;
        RECT 28.8 9.06 28.9 9.16 ;
        RECT 28.8 8.83 28.9 8.93 ;
        RECT 28.8 8.6 28.9 8.7 ;
        RECT 28.8 8.37 28.9 8.47 ;
        RECT 28.8 8.14 28.9 8.24 ;
        RECT 28.8 7.91 28.9 8.01 ;
        RECT 28.8 7.68 28.9 7.78 ;
        RECT 28.8 7.45 28.9 7.55 ;
        RECT 28.8 7.22 28.9 7.32 ;
        RECT 28.8 0.8 28.9 0.9 ;
        RECT 28.8 0.445 28.9 0.545 ;
        RECT 28.8 -0.545 28.9 -0.445 ;
        RECT 28.8 -0.9 28.9 -0.8 ;
        RECT 28.8 -2.43 28.9 -2.33 ;
        RECT 28.8 -2.785 28.9 -2.685 ;
        RECT 28.8 -3.775 28.9 -3.675 ;
        RECT 28.8 -4.13 28.9 -4.03 ;
        RECT 28.8 -5.66 28.9 -5.56 ;
        RECT 28.8 -6.015 28.9 -5.915 ;
        RECT 28.8 -7.005 28.9 -6.905 ;
        RECT 28.8 -7.36 28.9 -7.26 ;
        RECT 28.8 -8.89 28.9 -8.79 ;
        RECT 28.8 -9.245 28.9 -9.145 ;
        RECT 28.8 -10.235 28.9 -10.135 ;
        RECT 28.8 -10.59 28.9 -10.49 ;
        RECT 28.8 -12.12 28.9 -12.02 ;
        RECT 28.8 -12.475 28.9 -12.375 ;
        RECT 28.8 -13.465 28.9 -13.365 ;
        RECT 28.8 -13.82 28.9 -13.72 ;
        RECT 28.8 -15.35 28.9 -15.25 ;
        RECT 28.8 -15.705 28.9 -15.605 ;
        RECT 28.8 -16.695 28.9 -16.595 ;
        RECT 28.8 -17.05 28.9 -16.95 ;
        RECT 28.8 -18.58 28.9 -18.48 ;
        RECT 28.8 -18.935 28.9 -18.835 ;
        RECT 28.8 -19.925 28.9 -19.825 ;
        RECT 28.8 -20.28 28.9 -20.18 ;
        RECT 28.8 -21.81 28.9 -21.71 ;
        RECT 28.8 -22.165 28.9 -22.065 ;
        RECT 28.8 -23.155 28.9 -23.055 ;
        RECT 28.8 -23.51 28.9 -23.41 ;
        RECT 28.8 -25.04 28.9 -24.94 ;
        RECT 28.8 -25.395 28.9 -25.295 ;
        RECT 28.8 -26.385 28.9 -26.285 ;
        RECT 28.8 -26.74 28.9 -26.64 ;
        RECT 28.8 -28.27 28.9 -28.17 ;
        RECT 28.8 -28.625 28.9 -28.525 ;
        RECT 28.8 -29.615 28.9 -29.515 ;
        RECT 28.8 -29.97 28.9 -29.87 ;
        RECT 28.8 -31.5 28.9 -31.4 ;
        RECT 28.8 -31.855 28.9 -31.755 ;
        RECT 28.8 -32.845 28.9 -32.745 ;
        RECT 28.8 -33.2 28.9 -33.1 ;
        RECT 28.8 -34.73 28.9 -34.63 ;
        RECT 28.8 -35.085 28.9 -34.985 ;
        RECT 28.8 -36.075 28.9 -35.975 ;
        RECT 28.8 -36.43 28.9 -36.33 ;
        RECT 28.8 -37.96 28.9 -37.86 ;
        RECT 28.8 -38.315 28.9 -38.215 ;
        RECT 28.8 -39.305 28.9 -39.205 ;
        RECT 28.8 -39.66 28.9 -39.56 ;
        RECT 28.8 -41.19 28.9 -41.09 ;
        RECT 28.8 -41.545 28.9 -41.445 ;
        RECT 28.8 -42.535 28.9 -42.435 ;
        RECT 28.8 -42.89 28.9 -42.79 ;
        RECT 28.8 -44.42 28.9 -44.32 ;
        RECT 28.8 -44.775 28.9 -44.675 ;
        RECT 28.8 -45.765 28.9 -45.665 ;
        RECT 28.8 -46.12 28.9 -46.02 ;
        RECT 28.8 -47.65 28.9 -47.55 ;
        RECT 28.8 -48.005 28.9 -47.905 ;
        RECT 28.8 -48.995 28.9 -48.895 ;
        RECT 28.8 -49.35 28.9 -49.25 ;
        RECT 30 9.75 30.1 9.85 ;
        RECT 30 9.52 30.1 9.62 ;
        RECT 30 9.29 30.1 9.39 ;
        RECT 30 9.06 30.1 9.16 ;
        RECT 30 8.83 30.1 8.93 ;
        RECT 30 8.6 30.1 8.7 ;
        RECT 30 8.37 30.1 8.47 ;
        RECT 30 8.14 30.1 8.24 ;
        RECT 30 7.91 30.1 8.01 ;
        RECT 30 7.68 30.1 7.78 ;
        RECT 30 7.45 30.1 7.55 ;
        RECT 30 7.22 30.1 7.32 ;
        RECT 30 0.8 30.1 0.9 ;
        RECT 30 0.445 30.1 0.545 ;
        RECT 30 -0.545 30.1 -0.445 ;
        RECT 30 -0.9 30.1 -0.8 ;
        RECT 30 -2.43 30.1 -2.33 ;
        RECT 30 -2.785 30.1 -2.685 ;
        RECT 30 -3.775 30.1 -3.675 ;
        RECT 30 -4.13 30.1 -4.03 ;
        RECT 30 -5.66 30.1 -5.56 ;
        RECT 30 -6.015 30.1 -5.915 ;
        RECT 30 -7.005 30.1 -6.905 ;
        RECT 30 -7.36 30.1 -7.26 ;
        RECT 30 -8.89 30.1 -8.79 ;
        RECT 30 -9.245 30.1 -9.145 ;
        RECT 30 -10.235 30.1 -10.135 ;
        RECT 30 -10.59 30.1 -10.49 ;
        RECT 30 -12.12 30.1 -12.02 ;
        RECT 30 -12.475 30.1 -12.375 ;
        RECT 30 -13.465 30.1 -13.365 ;
        RECT 30 -13.82 30.1 -13.72 ;
        RECT 30 -15.35 30.1 -15.25 ;
        RECT 30 -15.705 30.1 -15.605 ;
        RECT 30 -16.695 30.1 -16.595 ;
        RECT 30 -17.05 30.1 -16.95 ;
        RECT 30 -18.58 30.1 -18.48 ;
        RECT 30 -18.935 30.1 -18.835 ;
        RECT 30 -19.925 30.1 -19.825 ;
        RECT 30 -20.28 30.1 -20.18 ;
        RECT 30 -21.81 30.1 -21.71 ;
        RECT 30 -22.165 30.1 -22.065 ;
        RECT 30 -23.155 30.1 -23.055 ;
        RECT 30 -23.51 30.1 -23.41 ;
        RECT 30 -25.04 30.1 -24.94 ;
        RECT 30 -25.395 30.1 -25.295 ;
        RECT 30 -26.385 30.1 -26.285 ;
        RECT 30 -26.74 30.1 -26.64 ;
        RECT 30 -28.27 30.1 -28.17 ;
        RECT 30 -28.625 30.1 -28.525 ;
        RECT 30 -29.615 30.1 -29.515 ;
        RECT 30 -29.97 30.1 -29.87 ;
        RECT 30 -31.5 30.1 -31.4 ;
        RECT 30 -31.855 30.1 -31.755 ;
        RECT 30 -32.845 30.1 -32.745 ;
        RECT 30 -33.2 30.1 -33.1 ;
        RECT 30 -34.73 30.1 -34.63 ;
        RECT 30 -35.085 30.1 -34.985 ;
        RECT 30 -36.075 30.1 -35.975 ;
        RECT 30 -36.43 30.1 -36.33 ;
        RECT 30 -37.96 30.1 -37.86 ;
        RECT 30 -38.315 30.1 -38.215 ;
        RECT 30 -39.305 30.1 -39.205 ;
        RECT 30 -39.66 30.1 -39.56 ;
        RECT 30 -41.19 30.1 -41.09 ;
        RECT 30 -41.545 30.1 -41.445 ;
        RECT 30 -42.535 30.1 -42.435 ;
        RECT 30 -42.89 30.1 -42.79 ;
        RECT 30 -44.42 30.1 -44.32 ;
        RECT 30 -44.775 30.1 -44.675 ;
        RECT 30 -45.765 30.1 -45.665 ;
        RECT 30 -46.12 30.1 -46.02 ;
        RECT 30 -47.65 30.1 -47.55 ;
        RECT 30 -48.005 30.1 -47.905 ;
        RECT 30 -48.995 30.1 -48.895 ;
        RECT 30 -49.35 30.1 -49.25 ;
        RECT 31.2 9.75 31.3 9.85 ;
        RECT 31.2 9.52 31.3 9.62 ;
        RECT 31.2 9.29 31.3 9.39 ;
        RECT 31.2 9.06 31.3 9.16 ;
        RECT 31.2 8.83 31.3 8.93 ;
        RECT 31.2 8.6 31.3 8.7 ;
        RECT 31.2 8.37 31.3 8.47 ;
        RECT 31.2 8.14 31.3 8.24 ;
        RECT 31.2 7.91 31.3 8.01 ;
        RECT 31.2 7.68 31.3 7.78 ;
        RECT 31.2 7.45 31.3 7.55 ;
        RECT 31.2 7.22 31.3 7.32 ;
        RECT 31.2 0.8 31.3 0.9 ;
        RECT 31.2 0.445 31.3 0.545 ;
        RECT 31.2 -0.545 31.3 -0.445 ;
        RECT 31.2 -0.9 31.3 -0.8 ;
        RECT 31.2 -2.43 31.3 -2.33 ;
        RECT 31.2 -2.785 31.3 -2.685 ;
        RECT 31.2 -3.775 31.3 -3.675 ;
        RECT 31.2 -4.13 31.3 -4.03 ;
        RECT 31.2 -5.66 31.3 -5.56 ;
        RECT 31.2 -6.015 31.3 -5.915 ;
        RECT 31.2 -7.005 31.3 -6.905 ;
        RECT 31.2 -7.36 31.3 -7.26 ;
        RECT 31.2 -8.89 31.3 -8.79 ;
        RECT 31.2 -9.245 31.3 -9.145 ;
        RECT 31.2 -10.235 31.3 -10.135 ;
        RECT 31.2 -10.59 31.3 -10.49 ;
        RECT 31.2 -12.12 31.3 -12.02 ;
        RECT 31.2 -12.475 31.3 -12.375 ;
        RECT 31.2 -13.465 31.3 -13.365 ;
        RECT 31.2 -13.82 31.3 -13.72 ;
        RECT 31.2 -15.35 31.3 -15.25 ;
        RECT 31.2 -15.705 31.3 -15.605 ;
        RECT 31.2 -16.695 31.3 -16.595 ;
        RECT 31.2 -17.05 31.3 -16.95 ;
        RECT 31.2 -18.58 31.3 -18.48 ;
        RECT 31.2 -18.935 31.3 -18.835 ;
        RECT 31.2 -19.925 31.3 -19.825 ;
        RECT 31.2 -20.28 31.3 -20.18 ;
        RECT 31.2 -21.81 31.3 -21.71 ;
        RECT 31.2 -22.165 31.3 -22.065 ;
        RECT 31.2 -23.155 31.3 -23.055 ;
        RECT 31.2 -23.51 31.3 -23.41 ;
        RECT 31.2 -25.04 31.3 -24.94 ;
        RECT 31.2 -25.395 31.3 -25.295 ;
        RECT 31.2 -26.385 31.3 -26.285 ;
        RECT 31.2 -26.74 31.3 -26.64 ;
        RECT 31.2 -28.27 31.3 -28.17 ;
        RECT 31.2 -28.625 31.3 -28.525 ;
        RECT 31.2 -29.615 31.3 -29.515 ;
        RECT 31.2 -29.97 31.3 -29.87 ;
        RECT 31.2 -31.5 31.3 -31.4 ;
        RECT 31.2 -31.855 31.3 -31.755 ;
        RECT 31.2 -32.845 31.3 -32.745 ;
        RECT 31.2 -33.2 31.3 -33.1 ;
        RECT 31.2 -34.73 31.3 -34.63 ;
        RECT 31.2 -35.085 31.3 -34.985 ;
        RECT 31.2 -36.075 31.3 -35.975 ;
        RECT 31.2 -36.43 31.3 -36.33 ;
        RECT 31.2 -37.96 31.3 -37.86 ;
        RECT 31.2 -38.315 31.3 -38.215 ;
        RECT 31.2 -39.305 31.3 -39.205 ;
        RECT 31.2 -39.66 31.3 -39.56 ;
        RECT 31.2 -41.19 31.3 -41.09 ;
        RECT 31.2 -41.545 31.3 -41.445 ;
        RECT 31.2 -42.535 31.3 -42.435 ;
        RECT 31.2 -42.89 31.3 -42.79 ;
        RECT 31.2 -44.42 31.3 -44.32 ;
        RECT 31.2 -44.775 31.3 -44.675 ;
        RECT 31.2 -45.765 31.3 -45.665 ;
        RECT 31.2 -46.12 31.3 -46.02 ;
        RECT 31.2 -47.65 31.3 -47.55 ;
        RECT 31.2 -48.005 31.3 -47.905 ;
        RECT 31.2 -48.995 31.3 -48.895 ;
        RECT 31.2 -49.35 31.3 -49.25 ;
        RECT 32.4 9.75 32.5 9.85 ;
        RECT 32.4 9.52 32.5 9.62 ;
        RECT 32.4 9.29 32.5 9.39 ;
        RECT 32.4 9.06 32.5 9.16 ;
        RECT 32.4 8.83 32.5 8.93 ;
        RECT 32.4 8.6 32.5 8.7 ;
        RECT 32.4 8.37 32.5 8.47 ;
        RECT 32.4 8.14 32.5 8.24 ;
        RECT 32.4 7.91 32.5 8.01 ;
        RECT 32.4 7.68 32.5 7.78 ;
        RECT 32.4 7.45 32.5 7.55 ;
        RECT 32.4 7.22 32.5 7.32 ;
        RECT 32.4 0.8 32.5 0.9 ;
        RECT 32.4 0.445 32.5 0.545 ;
        RECT 32.4 -0.545 32.5 -0.445 ;
        RECT 32.4 -0.9 32.5 -0.8 ;
        RECT 32.4 -2.43 32.5 -2.33 ;
        RECT 32.4 -2.785 32.5 -2.685 ;
        RECT 32.4 -3.775 32.5 -3.675 ;
        RECT 32.4 -4.13 32.5 -4.03 ;
        RECT 32.4 -5.66 32.5 -5.56 ;
        RECT 32.4 -6.015 32.5 -5.915 ;
        RECT 32.4 -7.005 32.5 -6.905 ;
        RECT 32.4 -7.36 32.5 -7.26 ;
        RECT 32.4 -8.89 32.5 -8.79 ;
        RECT 32.4 -9.245 32.5 -9.145 ;
        RECT 32.4 -10.235 32.5 -10.135 ;
        RECT 32.4 -10.59 32.5 -10.49 ;
        RECT 32.4 -12.12 32.5 -12.02 ;
        RECT 32.4 -12.475 32.5 -12.375 ;
        RECT 32.4 -13.465 32.5 -13.365 ;
        RECT 32.4 -13.82 32.5 -13.72 ;
        RECT 32.4 -15.35 32.5 -15.25 ;
        RECT 32.4 -15.705 32.5 -15.605 ;
        RECT 32.4 -16.695 32.5 -16.595 ;
        RECT 32.4 -17.05 32.5 -16.95 ;
        RECT 32.4 -18.58 32.5 -18.48 ;
        RECT 32.4 -18.935 32.5 -18.835 ;
        RECT 32.4 -19.925 32.5 -19.825 ;
        RECT 32.4 -20.28 32.5 -20.18 ;
        RECT 32.4 -21.81 32.5 -21.71 ;
        RECT 32.4 -22.165 32.5 -22.065 ;
        RECT 32.4 -23.155 32.5 -23.055 ;
        RECT 32.4 -23.51 32.5 -23.41 ;
        RECT 32.4 -25.04 32.5 -24.94 ;
        RECT 32.4 -25.395 32.5 -25.295 ;
        RECT 32.4 -26.385 32.5 -26.285 ;
        RECT 32.4 -26.74 32.5 -26.64 ;
        RECT 32.4 -28.27 32.5 -28.17 ;
        RECT 32.4 -28.625 32.5 -28.525 ;
        RECT 32.4 -29.615 32.5 -29.515 ;
        RECT 32.4 -29.97 32.5 -29.87 ;
        RECT 32.4 -31.5 32.5 -31.4 ;
        RECT 32.4 -31.855 32.5 -31.755 ;
        RECT 32.4 -32.845 32.5 -32.745 ;
        RECT 32.4 -33.2 32.5 -33.1 ;
        RECT 32.4 -34.73 32.5 -34.63 ;
        RECT 32.4 -35.085 32.5 -34.985 ;
        RECT 32.4 -36.075 32.5 -35.975 ;
        RECT 32.4 -36.43 32.5 -36.33 ;
        RECT 32.4 -37.96 32.5 -37.86 ;
        RECT 32.4 -38.315 32.5 -38.215 ;
        RECT 32.4 -39.305 32.5 -39.205 ;
        RECT 32.4 -39.66 32.5 -39.56 ;
        RECT 32.4 -41.19 32.5 -41.09 ;
        RECT 32.4 -41.545 32.5 -41.445 ;
        RECT 32.4 -42.535 32.5 -42.435 ;
        RECT 32.4 -42.89 32.5 -42.79 ;
        RECT 32.4 -44.42 32.5 -44.32 ;
        RECT 32.4 -44.775 32.5 -44.675 ;
        RECT 32.4 -45.765 32.5 -45.665 ;
        RECT 32.4 -46.12 32.5 -46.02 ;
        RECT 32.4 -47.65 32.5 -47.55 ;
        RECT 32.4 -48.005 32.5 -47.905 ;
        RECT 32.4 -48.995 32.5 -48.895 ;
        RECT 32.4 -49.35 32.5 -49.25 ;
        RECT 33.6 9.75 33.7 9.85 ;
        RECT 33.6 9.52 33.7 9.62 ;
        RECT 33.6 9.29 33.7 9.39 ;
        RECT 33.6 9.06 33.7 9.16 ;
        RECT 33.6 8.83 33.7 8.93 ;
        RECT 33.6 8.6 33.7 8.7 ;
        RECT 33.6 8.37 33.7 8.47 ;
        RECT 33.6 8.14 33.7 8.24 ;
        RECT 33.6 7.91 33.7 8.01 ;
        RECT 33.6 7.68 33.7 7.78 ;
        RECT 33.6 7.45 33.7 7.55 ;
        RECT 33.6 7.22 33.7 7.32 ;
        RECT 33.6 0.8 33.7 0.9 ;
        RECT 33.6 0.445 33.7 0.545 ;
        RECT 33.6 -0.545 33.7 -0.445 ;
        RECT 33.6 -0.9 33.7 -0.8 ;
        RECT 33.6 -2.43 33.7 -2.33 ;
        RECT 33.6 -2.785 33.7 -2.685 ;
        RECT 33.6 -3.775 33.7 -3.675 ;
        RECT 33.6 -4.13 33.7 -4.03 ;
        RECT 33.6 -5.66 33.7 -5.56 ;
        RECT 33.6 -6.015 33.7 -5.915 ;
        RECT 33.6 -7.005 33.7 -6.905 ;
        RECT 33.6 -7.36 33.7 -7.26 ;
        RECT 33.6 -8.89 33.7 -8.79 ;
        RECT 33.6 -9.245 33.7 -9.145 ;
        RECT 33.6 -10.235 33.7 -10.135 ;
        RECT 33.6 -10.59 33.7 -10.49 ;
        RECT 33.6 -12.12 33.7 -12.02 ;
        RECT 33.6 -12.475 33.7 -12.375 ;
        RECT 33.6 -13.465 33.7 -13.365 ;
        RECT 33.6 -13.82 33.7 -13.72 ;
        RECT 33.6 -15.35 33.7 -15.25 ;
        RECT 33.6 -15.705 33.7 -15.605 ;
        RECT 33.6 -16.695 33.7 -16.595 ;
        RECT 33.6 -17.05 33.7 -16.95 ;
        RECT 33.6 -18.58 33.7 -18.48 ;
        RECT 33.6 -18.935 33.7 -18.835 ;
        RECT 33.6 -19.925 33.7 -19.825 ;
        RECT 33.6 -20.28 33.7 -20.18 ;
        RECT 33.6 -21.81 33.7 -21.71 ;
        RECT 33.6 -22.165 33.7 -22.065 ;
        RECT 33.6 -23.155 33.7 -23.055 ;
        RECT 33.6 -23.51 33.7 -23.41 ;
        RECT 33.6 -25.04 33.7 -24.94 ;
        RECT 33.6 -25.395 33.7 -25.295 ;
        RECT 33.6 -26.385 33.7 -26.285 ;
        RECT 33.6 -26.74 33.7 -26.64 ;
        RECT 33.6 -28.27 33.7 -28.17 ;
        RECT 33.6 -28.625 33.7 -28.525 ;
        RECT 33.6 -29.615 33.7 -29.515 ;
        RECT 33.6 -29.97 33.7 -29.87 ;
        RECT 33.6 -31.5 33.7 -31.4 ;
        RECT 33.6 -31.855 33.7 -31.755 ;
        RECT 33.6 -32.845 33.7 -32.745 ;
        RECT 33.6 -33.2 33.7 -33.1 ;
        RECT 33.6 -34.73 33.7 -34.63 ;
        RECT 33.6 -35.085 33.7 -34.985 ;
        RECT 33.6 -36.075 33.7 -35.975 ;
        RECT 33.6 -36.43 33.7 -36.33 ;
        RECT 33.6 -37.96 33.7 -37.86 ;
        RECT 33.6 -38.315 33.7 -38.215 ;
        RECT 33.6 -39.305 33.7 -39.205 ;
        RECT 33.6 -39.66 33.7 -39.56 ;
        RECT 33.6 -41.19 33.7 -41.09 ;
        RECT 33.6 -41.545 33.7 -41.445 ;
        RECT 33.6 -42.535 33.7 -42.435 ;
        RECT 33.6 -42.89 33.7 -42.79 ;
        RECT 33.6 -44.42 33.7 -44.32 ;
        RECT 33.6 -44.775 33.7 -44.675 ;
        RECT 33.6 -45.765 33.7 -45.665 ;
        RECT 33.6 -46.12 33.7 -46.02 ;
        RECT 33.6 -47.65 33.7 -47.55 ;
        RECT 33.6 -48.005 33.7 -47.905 ;
        RECT 33.6 -48.995 33.7 -48.895 ;
        RECT 33.6 -49.35 33.7 -49.25 ;
        RECT 34.8 9.75 34.9 9.85 ;
        RECT 34.8 9.52 34.9 9.62 ;
        RECT 34.8 9.29 34.9 9.39 ;
        RECT 34.8 9.06 34.9 9.16 ;
        RECT 34.8 8.83 34.9 8.93 ;
        RECT 34.8 8.6 34.9 8.7 ;
        RECT 34.8 8.37 34.9 8.47 ;
        RECT 34.8 8.14 34.9 8.24 ;
        RECT 34.8 7.91 34.9 8.01 ;
        RECT 34.8 7.68 34.9 7.78 ;
        RECT 34.8 7.45 34.9 7.55 ;
        RECT 34.8 7.22 34.9 7.32 ;
        RECT 34.8 0.8 34.9 0.9 ;
        RECT 34.8 0.445 34.9 0.545 ;
        RECT 34.8 -0.545 34.9 -0.445 ;
        RECT 34.8 -0.9 34.9 -0.8 ;
        RECT 34.8 -2.43 34.9 -2.33 ;
        RECT 34.8 -2.785 34.9 -2.685 ;
        RECT 34.8 -3.775 34.9 -3.675 ;
        RECT 34.8 -4.13 34.9 -4.03 ;
        RECT 34.8 -5.66 34.9 -5.56 ;
        RECT 34.8 -6.015 34.9 -5.915 ;
        RECT 34.8 -7.005 34.9 -6.905 ;
        RECT 34.8 -7.36 34.9 -7.26 ;
        RECT 34.8 -8.89 34.9 -8.79 ;
        RECT 34.8 -9.245 34.9 -9.145 ;
        RECT 34.8 -10.235 34.9 -10.135 ;
        RECT 34.8 -10.59 34.9 -10.49 ;
        RECT 34.8 -12.12 34.9 -12.02 ;
        RECT 34.8 -12.475 34.9 -12.375 ;
        RECT 34.8 -13.465 34.9 -13.365 ;
        RECT 34.8 -13.82 34.9 -13.72 ;
        RECT 34.8 -15.35 34.9 -15.25 ;
        RECT 34.8 -15.705 34.9 -15.605 ;
        RECT 34.8 -16.695 34.9 -16.595 ;
        RECT 34.8 -17.05 34.9 -16.95 ;
        RECT 34.8 -18.58 34.9 -18.48 ;
        RECT 34.8 -18.935 34.9 -18.835 ;
        RECT 34.8 -19.925 34.9 -19.825 ;
        RECT 34.8 -20.28 34.9 -20.18 ;
        RECT 34.8 -21.81 34.9 -21.71 ;
        RECT 34.8 -22.165 34.9 -22.065 ;
        RECT 34.8 -23.155 34.9 -23.055 ;
        RECT 34.8 -23.51 34.9 -23.41 ;
        RECT 34.8 -25.04 34.9 -24.94 ;
        RECT 34.8 -25.395 34.9 -25.295 ;
        RECT 34.8 -26.385 34.9 -26.285 ;
        RECT 34.8 -26.74 34.9 -26.64 ;
        RECT 34.8 -28.27 34.9 -28.17 ;
        RECT 34.8 -28.625 34.9 -28.525 ;
        RECT 34.8 -29.615 34.9 -29.515 ;
        RECT 34.8 -29.97 34.9 -29.87 ;
        RECT 34.8 -31.5 34.9 -31.4 ;
        RECT 34.8 -31.855 34.9 -31.755 ;
        RECT 34.8 -32.845 34.9 -32.745 ;
        RECT 34.8 -33.2 34.9 -33.1 ;
        RECT 34.8 -34.73 34.9 -34.63 ;
        RECT 34.8 -35.085 34.9 -34.985 ;
        RECT 34.8 -36.075 34.9 -35.975 ;
        RECT 34.8 -36.43 34.9 -36.33 ;
        RECT 34.8 -37.96 34.9 -37.86 ;
        RECT 34.8 -38.315 34.9 -38.215 ;
        RECT 34.8 -39.305 34.9 -39.205 ;
        RECT 34.8 -39.66 34.9 -39.56 ;
        RECT 34.8 -41.19 34.9 -41.09 ;
        RECT 34.8 -41.545 34.9 -41.445 ;
        RECT 34.8 -42.535 34.9 -42.435 ;
        RECT 34.8 -42.89 34.9 -42.79 ;
        RECT 34.8 -44.42 34.9 -44.32 ;
        RECT 34.8 -44.775 34.9 -44.675 ;
        RECT 34.8 -45.765 34.9 -45.665 ;
        RECT 34.8 -46.12 34.9 -46.02 ;
        RECT 34.8 -47.65 34.9 -47.55 ;
        RECT 34.8 -48.005 34.9 -47.905 ;
        RECT 34.8 -48.995 34.9 -48.895 ;
        RECT 34.8 -49.35 34.9 -49.25 ;
        RECT 36 9.75 36.1 9.85 ;
        RECT 36 9.52 36.1 9.62 ;
        RECT 36 9.29 36.1 9.39 ;
        RECT 36 9.06 36.1 9.16 ;
        RECT 36 8.83 36.1 8.93 ;
        RECT 36 8.6 36.1 8.7 ;
        RECT 36 8.37 36.1 8.47 ;
        RECT 36 8.14 36.1 8.24 ;
        RECT 36 7.91 36.1 8.01 ;
        RECT 36 7.68 36.1 7.78 ;
        RECT 36 7.45 36.1 7.55 ;
        RECT 36 7.22 36.1 7.32 ;
        RECT 36 0.8 36.1 0.9 ;
        RECT 36 0.445 36.1 0.545 ;
        RECT 36 -0.545 36.1 -0.445 ;
        RECT 36 -0.9 36.1 -0.8 ;
        RECT 36 -2.43 36.1 -2.33 ;
        RECT 36 -2.785 36.1 -2.685 ;
        RECT 36 -3.775 36.1 -3.675 ;
        RECT 36 -4.13 36.1 -4.03 ;
        RECT 36 -5.66 36.1 -5.56 ;
        RECT 36 -6.015 36.1 -5.915 ;
        RECT 36 -7.005 36.1 -6.905 ;
        RECT 36 -7.36 36.1 -7.26 ;
        RECT 36 -8.89 36.1 -8.79 ;
        RECT 36 -9.245 36.1 -9.145 ;
        RECT 36 -10.235 36.1 -10.135 ;
        RECT 36 -10.59 36.1 -10.49 ;
        RECT 36 -12.12 36.1 -12.02 ;
        RECT 36 -12.475 36.1 -12.375 ;
        RECT 36 -13.465 36.1 -13.365 ;
        RECT 36 -13.82 36.1 -13.72 ;
        RECT 36 -15.35 36.1 -15.25 ;
        RECT 36 -15.705 36.1 -15.605 ;
        RECT 36 -16.695 36.1 -16.595 ;
        RECT 36 -17.05 36.1 -16.95 ;
        RECT 36 -18.58 36.1 -18.48 ;
        RECT 36 -18.935 36.1 -18.835 ;
        RECT 36 -19.925 36.1 -19.825 ;
        RECT 36 -20.28 36.1 -20.18 ;
        RECT 36 -21.81 36.1 -21.71 ;
        RECT 36 -22.165 36.1 -22.065 ;
        RECT 36 -23.155 36.1 -23.055 ;
        RECT 36 -23.51 36.1 -23.41 ;
        RECT 36 -25.04 36.1 -24.94 ;
        RECT 36 -25.395 36.1 -25.295 ;
        RECT 36 -26.385 36.1 -26.285 ;
        RECT 36 -26.74 36.1 -26.64 ;
        RECT 36 -28.27 36.1 -28.17 ;
        RECT 36 -28.625 36.1 -28.525 ;
        RECT 36 -29.615 36.1 -29.515 ;
        RECT 36 -29.97 36.1 -29.87 ;
        RECT 36 -31.5 36.1 -31.4 ;
        RECT 36 -31.855 36.1 -31.755 ;
        RECT 36 -32.845 36.1 -32.745 ;
        RECT 36 -33.2 36.1 -33.1 ;
        RECT 36 -34.73 36.1 -34.63 ;
        RECT 36 -35.085 36.1 -34.985 ;
        RECT 36 -36.075 36.1 -35.975 ;
        RECT 36 -36.43 36.1 -36.33 ;
        RECT 36 -37.96 36.1 -37.86 ;
        RECT 36 -38.315 36.1 -38.215 ;
        RECT 36 -39.305 36.1 -39.205 ;
        RECT 36 -39.66 36.1 -39.56 ;
        RECT 36 -41.19 36.1 -41.09 ;
        RECT 36 -41.545 36.1 -41.445 ;
        RECT 36 -42.535 36.1 -42.435 ;
        RECT 36 -42.89 36.1 -42.79 ;
        RECT 36 -44.42 36.1 -44.32 ;
        RECT 36 -44.775 36.1 -44.675 ;
        RECT 36 -45.765 36.1 -45.665 ;
        RECT 36 -46.12 36.1 -46.02 ;
        RECT 36 -47.65 36.1 -47.55 ;
        RECT 36 -48.005 36.1 -47.905 ;
        RECT 36 -48.995 36.1 -48.895 ;
        RECT 36 -49.35 36.1 -49.25 ;
        RECT 37.2 9.75 37.3 9.85 ;
        RECT 37.2 9.52 37.3 9.62 ;
        RECT 37.2 9.29 37.3 9.39 ;
        RECT 37.2 9.06 37.3 9.16 ;
        RECT 37.2 8.83 37.3 8.93 ;
        RECT 37.2 8.6 37.3 8.7 ;
        RECT 37.2 8.37 37.3 8.47 ;
        RECT 37.2 8.14 37.3 8.24 ;
        RECT 37.2 7.91 37.3 8.01 ;
        RECT 37.2 7.68 37.3 7.78 ;
        RECT 37.2 7.45 37.3 7.55 ;
        RECT 37.2 7.22 37.3 7.32 ;
        RECT 37.2 0.8 37.3 0.9 ;
        RECT 37.2 0.445 37.3 0.545 ;
        RECT 37.2 -0.545 37.3 -0.445 ;
        RECT 37.2 -0.9 37.3 -0.8 ;
        RECT 37.2 -2.43 37.3 -2.33 ;
        RECT 37.2 -2.785 37.3 -2.685 ;
        RECT 37.2 -3.775 37.3 -3.675 ;
        RECT 37.2 -4.13 37.3 -4.03 ;
        RECT 37.2 -5.66 37.3 -5.56 ;
        RECT 37.2 -6.015 37.3 -5.915 ;
        RECT 37.2 -7.005 37.3 -6.905 ;
        RECT 37.2 -7.36 37.3 -7.26 ;
        RECT 37.2 -8.89 37.3 -8.79 ;
        RECT 37.2 -9.245 37.3 -9.145 ;
        RECT 37.2 -10.235 37.3 -10.135 ;
        RECT 37.2 -10.59 37.3 -10.49 ;
        RECT 37.2 -12.12 37.3 -12.02 ;
        RECT 37.2 -12.475 37.3 -12.375 ;
        RECT 37.2 -13.465 37.3 -13.365 ;
        RECT 37.2 -13.82 37.3 -13.72 ;
        RECT 37.2 -15.35 37.3 -15.25 ;
        RECT 37.2 -15.705 37.3 -15.605 ;
        RECT 37.2 -16.695 37.3 -16.595 ;
        RECT 37.2 -17.05 37.3 -16.95 ;
        RECT 37.2 -18.58 37.3 -18.48 ;
        RECT 37.2 -18.935 37.3 -18.835 ;
        RECT 37.2 -19.925 37.3 -19.825 ;
        RECT 37.2 -20.28 37.3 -20.18 ;
        RECT 37.2 -21.81 37.3 -21.71 ;
        RECT 37.2 -22.165 37.3 -22.065 ;
        RECT 37.2 -23.155 37.3 -23.055 ;
        RECT 37.2 -23.51 37.3 -23.41 ;
        RECT 37.2 -25.04 37.3 -24.94 ;
        RECT 37.2 -25.395 37.3 -25.295 ;
        RECT 37.2 -26.385 37.3 -26.285 ;
        RECT 37.2 -26.74 37.3 -26.64 ;
        RECT 37.2 -28.27 37.3 -28.17 ;
        RECT 37.2 -28.625 37.3 -28.525 ;
        RECT 37.2 -29.615 37.3 -29.515 ;
        RECT 37.2 -29.97 37.3 -29.87 ;
        RECT 37.2 -31.5 37.3 -31.4 ;
        RECT 37.2 -31.855 37.3 -31.755 ;
        RECT 37.2 -32.845 37.3 -32.745 ;
        RECT 37.2 -33.2 37.3 -33.1 ;
        RECT 37.2 -34.73 37.3 -34.63 ;
        RECT 37.2 -35.085 37.3 -34.985 ;
        RECT 37.2 -36.075 37.3 -35.975 ;
        RECT 37.2 -36.43 37.3 -36.33 ;
        RECT 37.2 -37.96 37.3 -37.86 ;
        RECT 37.2 -38.315 37.3 -38.215 ;
        RECT 37.2 -39.305 37.3 -39.205 ;
        RECT 37.2 -39.66 37.3 -39.56 ;
        RECT 37.2 -41.19 37.3 -41.09 ;
        RECT 37.2 -41.545 37.3 -41.445 ;
        RECT 37.2 -42.535 37.3 -42.435 ;
        RECT 37.2 -42.89 37.3 -42.79 ;
        RECT 37.2 -44.42 37.3 -44.32 ;
        RECT 37.2 -44.775 37.3 -44.675 ;
        RECT 37.2 -45.765 37.3 -45.665 ;
        RECT 37.2 -46.12 37.3 -46.02 ;
        RECT 37.2 -47.65 37.3 -47.55 ;
        RECT 37.2 -48.005 37.3 -47.905 ;
        RECT 37.2 -48.995 37.3 -48.895 ;
        RECT 37.2 -49.35 37.3 -49.25 ;
        RECT 38.4 9.75 38.5 9.85 ;
        RECT 38.4 9.52 38.5 9.62 ;
        RECT 38.4 9.29 38.5 9.39 ;
        RECT 38.4 9.06 38.5 9.16 ;
        RECT 38.4 8.83 38.5 8.93 ;
        RECT 38.4 8.6 38.5 8.7 ;
        RECT 38.4 8.37 38.5 8.47 ;
        RECT 38.4 8.14 38.5 8.24 ;
        RECT 38.4 7.91 38.5 8.01 ;
        RECT 38.4 7.68 38.5 7.78 ;
        RECT 38.4 7.45 38.5 7.55 ;
        RECT 38.4 7.22 38.5 7.32 ;
        RECT 38.4 0.8 38.5 0.9 ;
        RECT 38.4 0.445 38.5 0.545 ;
        RECT 38.4 -0.545 38.5 -0.445 ;
        RECT 38.4 -0.9 38.5 -0.8 ;
        RECT 38.4 -2.43 38.5 -2.33 ;
        RECT 38.4 -2.785 38.5 -2.685 ;
        RECT 38.4 -3.775 38.5 -3.675 ;
        RECT 38.4 -4.13 38.5 -4.03 ;
        RECT 38.4 -5.66 38.5 -5.56 ;
        RECT 38.4 -6.015 38.5 -5.915 ;
        RECT 38.4 -7.005 38.5 -6.905 ;
        RECT 38.4 -7.36 38.5 -7.26 ;
        RECT 38.4 -8.89 38.5 -8.79 ;
        RECT 38.4 -9.245 38.5 -9.145 ;
        RECT 38.4 -10.235 38.5 -10.135 ;
        RECT 38.4 -10.59 38.5 -10.49 ;
        RECT 38.4 -12.12 38.5 -12.02 ;
        RECT 38.4 -12.475 38.5 -12.375 ;
        RECT 38.4 -13.465 38.5 -13.365 ;
        RECT 38.4 -13.82 38.5 -13.72 ;
        RECT 38.4 -15.35 38.5 -15.25 ;
        RECT 38.4 -15.705 38.5 -15.605 ;
        RECT 38.4 -16.695 38.5 -16.595 ;
        RECT 38.4 -17.05 38.5 -16.95 ;
        RECT 38.4 -18.58 38.5 -18.48 ;
        RECT 38.4 -18.935 38.5 -18.835 ;
        RECT 38.4 -19.925 38.5 -19.825 ;
        RECT 38.4 -20.28 38.5 -20.18 ;
        RECT 38.4 -21.81 38.5 -21.71 ;
        RECT 38.4 -22.165 38.5 -22.065 ;
        RECT 38.4 -23.155 38.5 -23.055 ;
        RECT 38.4 -23.51 38.5 -23.41 ;
        RECT 38.4 -25.04 38.5 -24.94 ;
        RECT 38.4 -25.395 38.5 -25.295 ;
        RECT 38.4 -26.385 38.5 -26.285 ;
        RECT 38.4 -26.74 38.5 -26.64 ;
        RECT 38.4 -28.27 38.5 -28.17 ;
        RECT 38.4 -28.625 38.5 -28.525 ;
        RECT 38.4 -29.615 38.5 -29.515 ;
        RECT 38.4 -29.97 38.5 -29.87 ;
        RECT 38.4 -31.5 38.5 -31.4 ;
        RECT 38.4 -31.855 38.5 -31.755 ;
        RECT 38.4 -32.845 38.5 -32.745 ;
        RECT 38.4 -33.2 38.5 -33.1 ;
        RECT 38.4 -34.73 38.5 -34.63 ;
        RECT 38.4 -35.085 38.5 -34.985 ;
        RECT 38.4 -36.075 38.5 -35.975 ;
        RECT 38.4 -36.43 38.5 -36.33 ;
        RECT 38.4 -37.96 38.5 -37.86 ;
        RECT 38.4 -38.315 38.5 -38.215 ;
        RECT 38.4 -39.305 38.5 -39.205 ;
        RECT 38.4 -39.66 38.5 -39.56 ;
        RECT 38.4 -41.19 38.5 -41.09 ;
        RECT 38.4 -41.545 38.5 -41.445 ;
        RECT 38.4 -42.535 38.5 -42.435 ;
        RECT 38.4 -42.89 38.5 -42.79 ;
        RECT 38.4 -44.42 38.5 -44.32 ;
        RECT 38.4 -44.775 38.5 -44.675 ;
        RECT 38.4 -45.765 38.5 -45.665 ;
        RECT 38.4 -46.12 38.5 -46.02 ;
        RECT 38.4 -47.65 38.5 -47.55 ;
        RECT 38.4 -48.005 38.5 -47.905 ;
        RECT 38.4 -48.995 38.5 -48.895 ;
        RECT 38.4 -49.35 38.5 -49.25 ;
        RECT 42.37 9.75 42.47 9.85 ;
        RECT 42.37 9.52 42.47 9.62 ;
        RECT 42.37 9.29 42.47 9.39 ;
        RECT 42.37 9.06 42.47 9.16 ;
        RECT 42.37 8.83 42.47 8.93 ;
        RECT 42.37 8.6 42.47 8.7 ;
        RECT 42.37 8.37 42.47 8.47 ;
        RECT 42.37 8.14 42.47 8.24 ;
        RECT 42.37 7.91 42.47 8.01 ;
        RECT 42.37 7.68 42.47 7.78 ;
        RECT 42.37 7.45 42.47 7.55 ;
        RECT 42.37 7.22 42.47 7.32 ;
        RECT 42.37 -58.385 42.47 -58.285 ;
        RECT 42.37 -63.645 42.47 -63.545 ;
        RECT 42.6 9.75 42.7 9.85 ;
        RECT 42.6 9.52 42.7 9.62 ;
        RECT 42.6 9.29 42.7 9.39 ;
        RECT 42.6 9.06 42.7 9.16 ;
        RECT 42.6 8.83 42.7 8.93 ;
        RECT 42.6 8.6 42.7 8.7 ;
        RECT 42.6 8.37 42.7 8.47 ;
        RECT 42.6 8.14 42.7 8.24 ;
        RECT 42.6 7.91 42.7 8.01 ;
        RECT 42.6 7.68 42.7 7.78 ;
        RECT 42.6 7.45 42.7 7.55 ;
        RECT 42.6 7.22 42.7 7.32 ;
        RECT 42.6 -58.385 42.7 -58.285 ;
        RECT 42.6 -63.645 42.7 -63.545 ;
        RECT 42.83 9.75 42.93 9.85 ;
        RECT 42.83 9.52 42.93 9.62 ;
        RECT 42.83 9.29 42.93 9.39 ;
        RECT 42.83 9.06 42.93 9.16 ;
        RECT 42.83 8.83 42.93 8.93 ;
        RECT 42.83 8.6 42.93 8.7 ;
        RECT 42.83 8.37 42.93 8.47 ;
        RECT 42.83 8.14 42.93 8.24 ;
        RECT 42.83 7.91 42.93 8.01 ;
        RECT 42.83 7.68 42.93 7.78 ;
        RECT 42.83 7.45 42.93 7.55 ;
        RECT 42.83 7.22 42.93 7.32 ;
        RECT 42.83 -58.385 42.93 -58.285 ;
        RECT 42.83 -63.645 42.93 -63.545 ;
        RECT 43.06 9.75 43.16 9.85 ;
        RECT 43.06 9.52 43.16 9.62 ;
        RECT 43.06 9.29 43.16 9.39 ;
        RECT 43.06 9.06 43.16 9.16 ;
        RECT 43.06 8.83 43.16 8.93 ;
        RECT 43.06 8.6 43.16 8.7 ;
        RECT 43.06 8.37 43.16 8.47 ;
        RECT 43.06 8.14 43.16 8.24 ;
        RECT 43.06 7.91 43.16 8.01 ;
        RECT 43.06 7.68 43.16 7.78 ;
        RECT 43.06 7.45 43.16 7.55 ;
        RECT 43.06 7.22 43.16 7.32 ;
        RECT 43.06 -58.385 43.16 -58.285 ;
        RECT 43.06 -63.645 43.16 -63.545 ;
        RECT 12 -28.27 12.1 -28.17 ;
        RECT 12 -28.625 12.1 -28.525 ;
        RECT 12 -29.615 12.1 -29.515 ;
        RECT 12 -29.97 12.1 -29.87 ;
        RECT 12 -31.5 12.1 -31.4 ;
        RECT 12 -31.855 12.1 -31.755 ;
        RECT 12 -32.845 12.1 -32.745 ;
        RECT 12 -33.2 12.1 -33.1 ;
        RECT 12 -34.73 12.1 -34.63 ;
        RECT 12 -35.085 12.1 -34.985 ;
        RECT 12 -36.075 12.1 -35.975 ;
        RECT 12 -36.43 12.1 -36.33 ;
        RECT 12 -37.96 12.1 -37.86 ;
        RECT 12 -38.315 12.1 -38.215 ;
        RECT 12 -39.305 12.1 -39.205 ;
        RECT 12 -39.66 12.1 -39.56 ;
        RECT 12 -41.19 12.1 -41.09 ;
        RECT 12 -41.545 12.1 -41.445 ;
        RECT 12 -42.535 12.1 -42.435 ;
        RECT 12 -42.89 12.1 -42.79 ;
        RECT 12 -44.42 12.1 -44.32 ;
        RECT 12 -44.775 12.1 -44.675 ;
        RECT 12 -45.765 12.1 -45.665 ;
        RECT 12 -46.12 12.1 -46.02 ;
        RECT 12 -47.65 12.1 -47.55 ;
        RECT 12 -48.005 12.1 -47.905 ;
        RECT 12 -48.995 12.1 -48.895 ;
        RECT 12 -49.35 12.1 -49.25 ;
        RECT 13.2 9.75 13.3 9.85 ;
        RECT 13.2 9.52 13.3 9.62 ;
        RECT 13.2 9.29 13.3 9.39 ;
        RECT 13.2 9.06 13.3 9.16 ;
        RECT 13.2 8.83 13.3 8.93 ;
        RECT 13.2 8.6 13.3 8.7 ;
        RECT 13.2 8.37 13.3 8.47 ;
        RECT 13.2 8.14 13.3 8.24 ;
        RECT 13.2 7.91 13.3 8.01 ;
        RECT 13.2 7.68 13.3 7.78 ;
        RECT 13.2 7.45 13.3 7.55 ;
        RECT 13.2 7.22 13.3 7.32 ;
        RECT 13.2 0.8 13.3 0.9 ;
        RECT 13.2 0.445 13.3 0.545 ;
        RECT 13.2 -0.545 13.3 -0.445 ;
        RECT 13.2 -0.9 13.3 -0.8 ;
        RECT 13.2 -2.43 13.3 -2.33 ;
        RECT 13.2 -2.785 13.3 -2.685 ;
        RECT 13.2 -3.775 13.3 -3.675 ;
        RECT 13.2 -4.13 13.3 -4.03 ;
        RECT 13.2 -5.66 13.3 -5.56 ;
        RECT 13.2 -6.015 13.3 -5.915 ;
        RECT 13.2 -7.005 13.3 -6.905 ;
        RECT 13.2 -7.36 13.3 -7.26 ;
        RECT 13.2 -8.89 13.3 -8.79 ;
        RECT 13.2 -9.245 13.3 -9.145 ;
        RECT 13.2 -10.235 13.3 -10.135 ;
        RECT 13.2 -10.59 13.3 -10.49 ;
        RECT 13.2 -12.12 13.3 -12.02 ;
        RECT 13.2 -12.475 13.3 -12.375 ;
        RECT 13.2 -13.465 13.3 -13.365 ;
        RECT 13.2 -13.82 13.3 -13.72 ;
        RECT 13.2 -15.35 13.3 -15.25 ;
        RECT 13.2 -15.705 13.3 -15.605 ;
        RECT 13.2 -16.695 13.3 -16.595 ;
        RECT 13.2 -17.05 13.3 -16.95 ;
        RECT 13.2 -18.58 13.3 -18.48 ;
        RECT 13.2 -18.935 13.3 -18.835 ;
        RECT 13.2 -19.925 13.3 -19.825 ;
        RECT 13.2 -20.28 13.3 -20.18 ;
        RECT 13.2 -21.81 13.3 -21.71 ;
        RECT 13.2 -22.165 13.3 -22.065 ;
        RECT 13.2 -23.155 13.3 -23.055 ;
        RECT 13.2 -23.51 13.3 -23.41 ;
        RECT 13.2 -25.04 13.3 -24.94 ;
        RECT 13.2 -25.395 13.3 -25.295 ;
        RECT 13.2 -26.385 13.3 -26.285 ;
        RECT 13.2 -26.74 13.3 -26.64 ;
        RECT 13.2 -28.27 13.3 -28.17 ;
        RECT 13.2 -28.625 13.3 -28.525 ;
        RECT 13.2 -29.615 13.3 -29.515 ;
        RECT 13.2 -29.97 13.3 -29.87 ;
        RECT 13.2 -31.5 13.3 -31.4 ;
        RECT 13.2 -31.855 13.3 -31.755 ;
        RECT 13.2 -32.845 13.3 -32.745 ;
        RECT 13.2 -33.2 13.3 -33.1 ;
        RECT 13.2 -34.73 13.3 -34.63 ;
        RECT 13.2 -35.085 13.3 -34.985 ;
        RECT 13.2 -36.075 13.3 -35.975 ;
        RECT 13.2 -36.43 13.3 -36.33 ;
        RECT 13.2 -37.96 13.3 -37.86 ;
        RECT 13.2 -38.315 13.3 -38.215 ;
        RECT 13.2 -39.305 13.3 -39.205 ;
        RECT 13.2 -39.66 13.3 -39.56 ;
        RECT 13.2 -41.19 13.3 -41.09 ;
        RECT 13.2 -41.545 13.3 -41.445 ;
        RECT 13.2 -42.535 13.3 -42.435 ;
        RECT 13.2 -42.89 13.3 -42.79 ;
        RECT 13.2 -44.42 13.3 -44.32 ;
        RECT 13.2 -44.775 13.3 -44.675 ;
        RECT 13.2 -45.765 13.3 -45.665 ;
        RECT 13.2 -46.12 13.3 -46.02 ;
        RECT 13.2 -47.65 13.3 -47.55 ;
        RECT 13.2 -48.005 13.3 -47.905 ;
        RECT 13.2 -48.995 13.3 -48.895 ;
        RECT 13.2 -49.35 13.3 -49.25 ;
        RECT 14.4 9.75 14.5 9.85 ;
        RECT 14.4 9.52 14.5 9.62 ;
        RECT 14.4 9.29 14.5 9.39 ;
        RECT 14.4 9.06 14.5 9.16 ;
        RECT 14.4 8.83 14.5 8.93 ;
        RECT 14.4 8.6 14.5 8.7 ;
        RECT 14.4 8.37 14.5 8.47 ;
        RECT 14.4 8.14 14.5 8.24 ;
        RECT 14.4 7.91 14.5 8.01 ;
        RECT 14.4 7.68 14.5 7.78 ;
        RECT 14.4 7.45 14.5 7.55 ;
        RECT 14.4 7.22 14.5 7.32 ;
        RECT 14.4 0.8 14.5 0.9 ;
        RECT 14.4 0.445 14.5 0.545 ;
        RECT 14.4 -0.545 14.5 -0.445 ;
        RECT 14.4 -0.9 14.5 -0.8 ;
        RECT 14.4 -2.43 14.5 -2.33 ;
        RECT 14.4 -2.785 14.5 -2.685 ;
        RECT 14.4 -3.775 14.5 -3.675 ;
        RECT 14.4 -4.13 14.5 -4.03 ;
        RECT 14.4 -5.66 14.5 -5.56 ;
        RECT 14.4 -6.015 14.5 -5.915 ;
        RECT 14.4 -7.005 14.5 -6.905 ;
        RECT 14.4 -7.36 14.5 -7.26 ;
        RECT 14.4 -8.89 14.5 -8.79 ;
        RECT 14.4 -9.245 14.5 -9.145 ;
        RECT 14.4 -10.235 14.5 -10.135 ;
        RECT 14.4 -10.59 14.5 -10.49 ;
        RECT 14.4 -12.12 14.5 -12.02 ;
        RECT 14.4 -12.475 14.5 -12.375 ;
        RECT 14.4 -13.465 14.5 -13.365 ;
        RECT 14.4 -13.82 14.5 -13.72 ;
        RECT 14.4 -15.35 14.5 -15.25 ;
        RECT 14.4 -15.705 14.5 -15.605 ;
        RECT 14.4 -16.695 14.5 -16.595 ;
        RECT 14.4 -17.05 14.5 -16.95 ;
        RECT 14.4 -18.58 14.5 -18.48 ;
        RECT 14.4 -18.935 14.5 -18.835 ;
        RECT 14.4 -19.925 14.5 -19.825 ;
        RECT 14.4 -20.28 14.5 -20.18 ;
        RECT 14.4 -21.81 14.5 -21.71 ;
        RECT 14.4 -22.165 14.5 -22.065 ;
        RECT 14.4 -23.155 14.5 -23.055 ;
        RECT 14.4 -23.51 14.5 -23.41 ;
        RECT 14.4 -25.04 14.5 -24.94 ;
        RECT 14.4 -25.395 14.5 -25.295 ;
        RECT 14.4 -26.385 14.5 -26.285 ;
        RECT 14.4 -26.74 14.5 -26.64 ;
        RECT 14.4 -28.27 14.5 -28.17 ;
        RECT 14.4 -28.625 14.5 -28.525 ;
        RECT 14.4 -29.615 14.5 -29.515 ;
        RECT 14.4 -29.97 14.5 -29.87 ;
        RECT 14.4 -31.5 14.5 -31.4 ;
        RECT 14.4 -31.855 14.5 -31.755 ;
        RECT 14.4 -32.845 14.5 -32.745 ;
        RECT 14.4 -33.2 14.5 -33.1 ;
        RECT 14.4 -34.73 14.5 -34.63 ;
        RECT 14.4 -35.085 14.5 -34.985 ;
        RECT 14.4 -36.075 14.5 -35.975 ;
        RECT 14.4 -36.43 14.5 -36.33 ;
        RECT 14.4 -37.96 14.5 -37.86 ;
        RECT 14.4 -38.315 14.5 -38.215 ;
        RECT 14.4 -39.305 14.5 -39.205 ;
        RECT 14.4 -39.66 14.5 -39.56 ;
        RECT 14.4 -41.19 14.5 -41.09 ;
        RECT 14.4 -41.545 14.5 -41.445 ;
        RECT 14.4 -42.535 14.5 -42.435 ;
        RECT 14.4 -42.89 14.5 -42.79 ;
        RECT 14.4 -44.42 14.5 -44.32 ;
        RECT 14.4 -44.775 14.5 -44.675 ;
        RECT 14.4 -45.765 14.5 -45.665 ;
        RECT 14.4 -46.12 14.5 -46.02 ;
        RECT 14.4 -47.65 14.5 -47.55 ;
        RECT 14.4 -48.005 14.5 -47.905 ;
        RECT 14.4 -48.995 14.5 -48.895 ;
        RECT 14.4 -49.35 14.5 -49.25 ;
        RECT 15.6 9.75 15.7 9.85 ;
        RECT 15.6 9.52 15.7 9.62 ;
        RECT 15.6 9.29 15.7 9.39 ;
        RECT 15.6 9.06 15.7 9.16 ;
        RECT 15.6 8.83 15.7 8.93 ;
        RECT 15.6 8.6 15.7 8.7 ;
        RECT 15.6 8.37 15.7 8.47 ;
        RECT 15.6 8.14 15.7 8.24 ;
        RECT 15.6 7.91 15.7 8.01 ;
        RECT 15.6 7.68 15.7 7.78 ;
        RECT 15.6 7.45 15.7 7.55 ;
        RECT 15.6 7.22 15.7 7.32 ;
        RECT 15.6 0.8 15.7 0.9 ;
        RECT 15.6 0.445 15.7 0.545 ;
        RECT 15.6 -0.545 15.7 -0.445 ;
        RECT 15.6 -0.9 15.7 -0.8 ;
        RECT 15.6 -2.43 15.7 -2.33 ;
        RECT 15.6 -2.785 15.7 -2.685 ;
        RECT 15.6 -3.775 15.7 -3.675 ;
        RECT 15.6 -4.13 15.7 -4.03 ;
        RECT 15.6 -5.66 15.7 -5.56 ;
        RECT 15.6 -6.015 15.7 -5.915 ;
        RECT 15.6 -7.005 15.7 -6.905 ;
        RECT 15.6 -7.36 15.7 -7.26 ;
        RECT 15.6 -8.89 15.7 -8.79 ;
        RECT 15.6 -9.245 15.7 -9.145 ;
        RECT 15.6 -10.235 15.7 -10.135 ;
        RECT 15.6 -10.59 15.7 -10.49 ;
        RECT 15.6 -12.12 15.7 -12.02 ;
        RECT 15.6 -12.475 15.7 -12.375 ;
        RECT 15.6 -13.465 15.7 -13.365 ;
        RECT 15.6 -13.82 15.7 -13.72 ;
        RECT 15.6 -15.35 15.7 -15.25 ;
        RECT 15.6 -15.705 15.7 -15.605 ;
        RECT 15.6 -16.695 15.7 -16.595 ;
        RECT 15.6 -17.05 15.7 -16.95 ;
        RECT 15.6 -18.58 15.7 -18.48 ;
        RECT 15.6 -18.935 15.7 -18.835 ;
        RECT 15.6 -19.925 15.7 -19.825 ;
        RECT 15.6 -20.28 15.7 -20.18 ;
        RECT 15.6 -21.81 15.7 -21.71 ;
        RECT 15.6 -22.165 15.7 -22.065 ;
        RECT 15.6 -23.155 15.7 -23.055 ;
        RECT 15.6 -23.51 15.7 -23.41 ;
        RECT 15.6 -25.04 15.7 -24.94 ;
        RECT 15.6 -25.395 15.7 -25.295 ;
        RECT 15.6 -26.385 15.7 -26.285 ;
        RECT 15.6 -26.74 15.7 -26.64 ;
        RECT 15.6 -28.27 15.7 -28.17 ;
        RECT 15.6 -28.625 15.7 -28.525 ;
        RECT 15.6 -29.615 15.7 -29.515 ;
        RECT 15.6 -29.97 15.7 -29.87 ;
        RECT 15.6 -31.5 15.7 -31.4 ;
        RECT 15.6 -31.855 15.7 -31.755 ;
        RECT 15.6 -32.845 15.7 -32.745 ;
        RECT 15.6 -33.2 15.7 -33.1 ;
        RECT 15.6 -34.73 15.7 -34.63 ;
        RECT 15.6 -35.085 15.7 -34.985 ;
        RECT 15.6 -36.075 15.7 -35.975 ;
        RECT 15.6 -36.43 15.7 -36.33 ;
        RECT 15.6 -37.96 15.7 -37.86 ;
        RECT 15.6 -38.315 15.7 -38.215 ;
        RECT 15.6 -39.305 15.7 -39.205 ;
        RECT 15.6 -39.66 15.7 -39.56 ;
        RECT 15.6 -41.19 15.7 -41.09 ;
        RECT 15.6 -41.545 15.7 -41.445 ;
        RECT 15.6 -42.535 15.7 -42.435 ;
        RECT 15.6 -42.89 15.7 -42.79 ;
        RECT 15.6 -44.42 15.7 -44.32 ;
        RECT 15.6 -44.775 15.7 -44.675 ;
        RECT 15.6 -45.765 15.7 -45.665 ;
        RECT 15.6 -46.12 15.7 -46.02 ;
        RECT 15.6 -47.65 15.7 -47.55 ;
        RECT 15.6 -48.005 15.7 -47.905 ;
        RECT 15.6 -48.995 15.7 -48.895 ;
        RECT 15.6 -49.35 15.7 -49.25 ;
        RECT 16.8 9.75 16.9 9.85 ;
        RECT 16.8 9.52 16.9 9.62 ;
        RECT 16.8 9.29 16.9 9.39 ;
        RECT 16.8 9.06 16.9 9.16 ;
        RECT 16.8 8.83 16.9 8.93 ;
        RECT 16.8 8.6 16.9 8.7 ;
        RECT 16.8 8.37 16.9 8.47 ;
        RECT 16.8 8.14 16.9 8.24 ;
        RECT 16.8 7.91 16.9 8.01 ;
        RECT 16.8 7.68 16.9 7.78 ;
        RECT 16.8 7.45 16.9 7.55 ;
        RECT 16.8 7.22 16.9 7.32 ;
        RECT 16.8 0.8 16.9 0.9 ;
        RECT 16.8 0.445 16.9 0.545 ;
        RECT 16.8 -0.545 16.9 -0.445 ;
        RECT 16.8 -0.9 16.9 -0.8 ;
        RECT 16.8 -2.43 16.9 -2.33 ;
        RECT 16.8 -2.785 16.9 -2.685 ;
        RECT 16.8 -3.775 16.9 -3.675 ;
        RECT 16.8 -4.13 16.9 -4.03 ;
        RECT 16.8 -5.66 16.9 -5.56 ;
        RECT 16.8 -6.015 16.9 -5.915 ;
        RECT 16.8 -7.005 16.9 -6.905 ;
        RECT 16.8 -7.36 16.9 -7.26 ;
        RECT 16.8 -8.89 16.9 -8.79 ;
        RECT 16.8 -9.245 16.9 -9.145 ;
        RECT 16.8 -10.235 16.9 -10.135 ;
        RECT 16.8 -10.59 16.9 -10.49 ;
        RECT 16.8 -12.12 16.9 -12.02 ;
        RECT 16.8 -12.475 16.9 -12.375 ;
        RECT 16.8 -13.465 16.9 -13.365 ;
        RECT 16.8 -13.82 16.9 -13.72 ;
        RECT 16.8 -15.35 16.9 -15.25 ;
        RECT 16.8 -15.705 16.9 -15.605 ;
        RECT 16.8 -16.695 16.9 -16.595 ;
        RECT 16.8 -17.05 16.9 -16.95 ;
        RECT 16.8 -18.58 16.9 -18.48 ;
        RECT 16.8 -18.935 16.9 -18.835 ;
        RECT 16.8 -19.925 16.9 -19.825 ;
        RECT 16.8 -20.28 16.9 -20.18 ;
        RECT 16.8 -21.81 16.9 -21.71 ;
        RECT 16.8 -22.165 16.9 -22.065 ;
        RECT 16.8 -23.155 16.9 -23.055 ;
        RECT 16.8 -23.51 16.9 -23.41 ;
        RECT 16.8 -25.04 16.9 -24.94 ;
        RECT 16.8 -25.395 16.9 -25.295 ;
        RECT 16.8 -26.385 16.9 -26.285 ;
        RECT 16.8 -26.74 16.9 -26.64 ;
        RECT 16.8 -28.27 16.9 -28.17 ;
        RECT 16.8 -28.625 16.9 -28.525 ;
        RECT 16.8 -29.615 16.9 -29.515 ;
        RECT 16.8 -29.97 16.9 -29.87 ;
        RECT 16.8 -31.5 16.9 -31.4 ;
        RECT 16.8 -31.855 16.9 -31.755 ;
        RECT 16.8 -32.845 16.9 -32.745 ;
        RECT 16.8 -33.2 16.9 -33.1 ;
        RECT 16.8 -34.73 16.9 -34.63 ;
        RECT 16.8 -35.085 16.9 -34.985 ;
        RECT 16.8 -36.075 16.9 -35.975 ;
        RECT 16.8 -36.43 16.9 -36.33 ;
        RECT 16.8 -37.96 16.9 -37.86 ;
        RECT 16.8 -38.315 16.9 -38.215 ;
        RECT 16.8 -39.305 16.9 -39.205 ;
        RECT 16.8 -39.66 16.9 -39.56 ;
        RECT 16.8 -41.19 16.9 -41.09 ;
        RECT 16.8 -41.545 16.9 -41.445 ;
        RECT 16.8 -42.535 16.9 -42.435 ;
        RECT 16.8 -42.89 16.9 -42.79 ;
        RECT 16.8 -44.42 16.9 -44.32 ;
        RECT 16.8 -44.775 16.9 -44.675 ;
        RECT 16.8 -45.765 16.9 -45.665 ;
        RECT 16.8 -46.12 16.9 -46.02 ;
        RECT 16.8 -47.65 16.9 -47.55 ;
        RECT 16.8 -48.005 16.9 -47.905 ;
        RECT 16.8 -48.995 16.9 -48.895 ;
        RECT 16.8 -49.35 16.9 -49.25 ;
        RECT 18 9.75 18.1 9.85 ;
        RECT 18 9.52 18.1 9.62 ;
        RECT 18 9.29 18.1 9.39 ;
        RECT 18 9.06 18.1 9.16 ;
        RECT 18 8.83 18.1 8.93 ;
        RECT 18 8.6 18.1 8.7 ;
        RECT 18 8.37 18.1 8.47 ;
        RECT 18 8.14 18.1 8.24 ;
        RECT 18 7.91 18.1 8.01 ;
        RECT 18 7.68 18.1 7.78 ;
        RECT 18 7.45 18.1 7.55 ;
        RECT 18 7.22 18.1 7.32 ;
        RECT 18 0.8 18.1 0.9 ;
        RECT 18 0.445 18.1 0.545 ;
        RECT 18 -0.545 18.1 -0.445 ;
        RECT 18 -0.9 18.1 -0.8 ;
        RECT 18 -2.43 18.1 -2.33 ;
        RECT 18 -2.785 18.1 -2.685 ;
        RECT 18 -3.775 18.1 -3.675 ;
        RECT 18 -4.13 18.1 -4.03 ;
        RECT 18 -5.66 18.1 -5.56 ;
        RECT 18 -6.015 18.1 -5.915 ;
        RECT 18 -7.005 18.1 -6.905 ;
        RECT 18 -7.36 18.1 -7.26 ;
        RECT 18 -8.89 18.1 -8.79 ;
        RECT 18 -9.245 18.1 -9.145 ;
        RECT 18 -10.235 18.1 -10.135 ;
        RECT 18 -10.59 18.1 -10.49 ;
        RECT 18 -12.12 18.1 -12.02 ;
        RECT 18 -12.475 18.1 -12.375 ;
        RECT 18 -13.465 18.1 -13.365 ;
        RECT 18 -13.82 18.1 -13.72 ;
        RECT 18 -15.35 18.1 -15.25 ;
        RECT 18 -15.705 18.1 -15.605 ;
        RECT 18 -16.695 18.1 -16.595 ;
        RECT 18 -17.05 18.1 -16.95 ;
        RECT 18 -18.58 18.1 -18.48 ;
        RECT 18 -18.935 18.1 -18.835 ;
        RECT 18 -19.925 18.1 -19.825 ;
        RECT 18 -20.28 18.1 -20.18 ;
        RECT 18 -21.81 18.1 -21.71 ;
        RECT 18 -22.165 18.1 -22.065 ;
        RECT 18 -23.155 18.1 -23.055 ;
        RECT 18 -23.51 18.1 -23.41 ;
        RECT 18 -25.04 18.1 -24.94 ;
        RECT 18 -25.395 18.1 -25.295 ;
        RECT 18 -26.385 18.1 -26.285 ;
        RECT 18 -26.74 18.1 -26.64 ;
        RECT 18 -28.27 18.1 -28.17 ;
        RECT 18 -28.625 18.1 -28.525 ;
        RECT 18 -29.615 18.1 -29.515 ;
        RECT 18 -29.97 18.1 -29.87 ;
        RECT 18 -31.5 18.1 -31.4 ;
        RECT 18 -31.855 18.1 -31.755 ;
        RECT 18 -32.845 18.1 -32.745 ;
        RECT 18 -33.2 18.1 -33.1 ;
        RECT 18 -34.73 18.1 -34.63 ;
        RECT 18 -35.085 18.1 -34.985 ;
        RECT 18 -36.075 18.1 -35.975 ;
        RECT 18 -36.43 18.1 -36.33 ;
        RECT 18 -37.96 18.1 -37.86 ;
        RECT 18 -38.315 18.1 -38.215 ;
        RECT 18 -39.305 18.1 -39.205 ;
        RECT 18 -39.66 18.1 -39.56 ;
        RECT 18 -41.19 18.1 -41.09 ;
        RECT 18 -41.545 18.1 -41.445 ;
        RECT 18 -42.535 18.1 -42.435 ;
        RECT 18 -42.89 18.1 -42.79 ;
        RECT 18 -44.42 18.1 -44.32 ;
        RECT 18 -44.775 18.1 -44.675 ;
        RECT 18 -45.765 18.1 -45.665 ;
        RECT 18 -46.12 18.1 -46.02 ;
        RECT 18 -47.65 18.1 -47.55 ;
        RECT 18 -48.005 18.1 -47.905 ;
        RECT 18 -48.995 18.1 -48.895 ;
        RECT 18 -49.35 18.1 -49.25 ;
        RECT 19.2 9.75 19.3 9.85 ;
        RECT 19.2 9.52 19.3 9.62 ;
        RECT 19.2 9.29 19.3 9.39 ;
        RECT 19.2 9.06 19.3 9.16 ;
        RECT 19.2 8.83 19.3 8.93 ;
        RECT 19.2 8.6 19.3 8.7 ;
        RECT 19.2 8.37 19.3 8.47 ;
        RECT 19.2 8.14 19.3 8.24 ;
        RECT 19.2 7.91 19.3 8.01 ;
        RECT 19.2 7.68 19.3 7.78 ;
        RECT 19.2 7.45 19.3 7.55 ;
        RECT 19.2 7.22 19.3 7.32 ;
        RECT 19.2 0.8 19.3 0.9 ;
        RECT 19.2 0.445 19.3 0.545 ;
        RECT 19.2 -0.545 19.3 -0.445 ;
        RECT 19.2 -0.9 19.3 -0.8 ;
        RECT 19.2 -2.43 19.3 -2.33 ;
        RECT 19.2 -2.785 19.3 -2.685 ;
        RECT 19.2 -3.775 19.3 -3.675 ;
        RECT 19.2 -4.13 19.3 -4.03 ;
        RECT 19.2 -5.66 19.3 -5.56 ;
        RECT 19.2 -6.015 19.3 -5.915 ;
        RECT 19.2 -7.005 19.3 -6.905 ;
        RECT 19.2 -7.36 19.3 -7.26 ;
        RECT 19.2 -8.89 19.3 -8.79 ;
        RECT 19.2 -9.245 19.3 -9.145 ;
        RECT 19.2 -10.235 19.3 -10.135 ;
        RECT 19.2 -10.59 19.3 -10.49 ;
        RECT 19.2 -12.12 19.3 -12.02 ;
        RECT 19.2 -12.475 19.3 -12.375 ;
        RECT 19.2 -13.465 19.3 -13.365 ;
        RECT 19.2 -13.82 19.3 -13.72 ;
        RECT 19.2 -15.35 19.3 -15.25 ;
        RECT 19.2 -15.705 19.3 -15.605 ;
        RECT 19.2 -16.695 19.3 -16.595 ;
        RECT 19.2 -17.05 19.3 -16.95 ;
        RECT 19.2 -18.58 19.3 -18.48 ;
        RECT 19.2 -18.935 19.3 -18.835 ;
        RECT 19.2 -19.925 19.3 -19.825 ;
        RECT 19.2 -20.28 19.3 -20.18 ;
        RECT 19.2 -21.81 19.3 -21.71 ;
        RECT 19.2 -22.165 19.3 -22.065 ;
        RECT 19.2 -23.155 19.3 -23.055 ;
        RECT 19.2 -23.51 19.3 -23.41 ;
        RECT 19.2 -25.04 19.3 -24.94 ;
        RECT 19.2 -25.395 19.3 -25.295 ;
        RECT 19.2 -26.385 19.3 -26.285 ;
        RECT 19.2 -26.74 19.3 -26.64 ;
        RECT 19.2 -28.27 19.3 -28.17 ;
        RECT 19.2 -28.625 19.3 -28.525 ;
        RECT 19.2 -29.615 19.3 -29.515 ;
        RECT 19.2 -29.97 19.3 -29.87 ;
        RECT 19.2 -31.5 19.3 -31.4 ;
        RECT 19.2 -31.855 19.3 -31.755 ;
        RECT 19.2 -32.845 19.3 -32.745 ;
        RECT 19.2 -33.2 19.3 -33.1 ;
        RECT 19.2 -34.73 19.3 -34.63 ;
        RECT 19.2 -35.085 19.3 -34.985 ;
        RECT 19.2 -36.075 19.3 -35.975 ;
        RECT 19.2 -36.43 19.3 -36.33 ;
        RECT 19.2 -37.96 19.3 -37.86 ;
        RECT 19.2 -38.315 19.3 -38.215 ;
        RECT 19.2 -39.305 19.3 -39.205 ;
        RECT 19.2 -39.66 19.3 -39.56 ;
        RECT 19.2 -41.19 19.3 -41.09 ;
        RECT 19.2 -41.545 19.3 -41.445 ;
        RECT 19.2 -42.535 19.3 -42.435 ;
        RECT 19.2 -42.89 19.3 -42.79 ;
        RECT 19.2 -44.42 19.3 -44.32 ;
        RECT 19.2 -44.775 19.3 -44.675 ;
        RECT 19.2 -45.765 19.3 -45.665 ;
        RECT 19.2 -46.12 19.3 -46.02 ;
        RECT 19.2 -47.65 19.3 -47.55 ;
        RECT 19.2 -48.005 19.3 -47.905 ;
        RECT 19.2 -48.995 19.3 -48.895 ;
        RECT 19.2 -49.35 19.3 -49.25 ;
        RECT 20.4 9.75 20.5 9.85 ;
        RECT 20.4 9.52 20.5 9.62 ;
        RECT 20.4 9.29 20.5 9.39 ;
        RECT 20.4 9.06 20.5 9.16 ;
        RECT 20.4 8.83 20.5 8.93 ;
        RECT 20.4 8.6 20.5 8.7 ;
        RECT 20.4 8.37 20.5 8.47 ;
        RECT 20.4 8.14 20.5 8.24 ;
        RECT 20.4 7.91 20.5 8.01 ;
        RECT 20.4 7.68 20.5 7.78 ;
        RECT 20.4 7.45 20.5 7.55 ;
        RECT 20.4 7.22 20.5 7.32 ;
        RECT 20.4 0.8 20.5 0.9 ;
        RECT 20.4 0.445 20.5 0.545 ;
        RECT 20.4 -0.545 20.5 -0.445 ;
        RECT 20.4 -0.9 20.5 -0.8 ;
        RECT 20.4 -2.43 20.5 -2.33 ;
        RECT 20.4 -2.785 20.5 -2.685 ;
        RECT 20.4 -3.775 20.5 -3.675 ;
        RECT 20.4 -4.13 20.5 -4.03 ;
        RECT 20.4 -5.66 20.5 -5.56 ;
        RECT 20.4 -6.015 20.5 -5.915 ;
        RECT 20.4 -7.005 20.5 -6.905 ;
        RECT 20.4 -7.36 20.5 -7.26 ;
        RECT 20.4 -8.89 20.5 -8.79 ;
        RECT 20.4 -9.245 20.5 -9.145 ;
        RECT 20.4 -10.235 20.5 -10.135 ;
        RECT 20.4 -10.59 20.5 -10.49 ;
        RECT 20.4 -12.12 20.5 -12.02 ;
        RECT 20.4 -12.475 20.5 -12.375 ;
        RECT 20.4 -13.465 20.5 -13.365 ;
        RECT 20.4 -13.82 20.5 -13.72 ;
        RECT 20.4 -15.35 20.5 -15.25 ;
        RECT 20.4 -15.705 20.5 -15.605 ;
        RECT 20.4 -16.695 20.5 -16.595 ;
        RECT 20.4 -17.05 20.5 -16.95 ;
        RECT 20.4 -18.58 20.5 -18.48 ;
        RECT 20.4 -18.935 20.5 -18.835 ;
        RECT 20.4 -19.925 20.5 -19.825 ;
        RECT 20.4 -20.28 20.5 -20.18 ;
        RECT 20.4 -21.81 20.5 -21.71 ;
        RECT 20.4 -22.165 20.5 -22.065 ;
        RECT 20.4 -23.155 20.5 -23.055 ;
        RECT 20.4 -23.51 20.5 -23.41 ;
        RECT 20.4 -25.04 20.5 -24.94 ;
        RECT 20.4 -25.395 20.5 -25.295 ;
        RECT 20.4 -26.385 20.5 -26.285 ;
        RECT 20.4 -26.74 20.5 -26.64 ;
        RECT 20.4 -28.27 20.5 -28.17 ;
        RECT 20.4 -28.625 20.5 -28.525 ;
        RECT 20.4 -29.615 20.5 -29.515 ;
        RECT 20.4 -29.97 20.5 -29.87 ;
        RECT 20.4 -31.5 20.5 -31.4 ;
        RECT 20.4 -31.855 20.5 -31.755 ;
        RECT 20.4 -32.845 20.5 -32.745 ;
        RECT 20.4 -33.2 20.5 -33.1 ;
        RECT 20.4 -34.73 20.5 -34.63 ;
        RECT 20.4 -35.085 20.5 -34.985 ;
        RECT 20.4 -36.075 20.5 -35.975 ;
        RECT 20.4 -36.43 20.5 -36.33 ;
        RECT 20.4 -37.96 20.5 -37.86 ;
        RECT 20.4 -38.315 20.5 -38.215 ;
        RECT 20.4 -39.305 20.5 -39.205 ;
        RECT 20.4 -39.66 20.5 -39.56 ;
        RECT 20.4 -41.19 20.5 -41.09 ;
        RECT 20.4 -41.545 20.5 -41.445 ;
        RECT 20.4 -42.535 20.5 -42.435 ;
        RECT 20.4 -42.89 20.5 -42.79 ;
        RECT 20.4 -44.42 20.5 -44.32 ;
        RECT 20.4 -44.775 20.5 -44.675 ;
        RECT 20.4 -45.765 20.5 -45.665 ;
        RECT 20.4 -46.12 20.5 -46.02 ;
        RECT 20.4 -47.65 20.5 -47.55 ;
        RECT 20.4 -48.005 20.5 -47.905 ;
        RECT 20.4 -48.995 20.5 -48.895 ;
        RECT 20.4 -49.35 20.5 -49.25 ;
        RECT 21.6 9.75 21.7 9.85 ;
        RECT 21.6 9.52 21.7 9.62 ;
        RECT 21.6 9.29 21.7 9.39 ;
        RECT 21.6 9.06 21.7 9.16 ;
        RECT 21.6 8.83 21.7 8.93 ;
        RECT 21.6 8.6 21.7 8.7 ;
        RECT 21.6 8.37 21.7 8.47 ;
        RECT 21.6 8.14 21.7 8.24 ;
        RECT 21.6 7.91 21.7 8.01 ;
        RECT 21.6 7.68 21.7 7.78 ;
        RECT 21.6 7.45 21.7 7.55 ;
        RECT 21.6 7.22 21.7 7.32 ;
        RECT 21.6 0.8 21.7 0.9 ;
        RECT 21.6 0.445 21.7 0.545 ;
        RECT 21.6 -0.545 21.7 -0.445 ;
        RECT 21.6 -0.9 21.7 -0.8 ;
        RECT 21.6 -2.43 21.7 -2.33 ;
        RECT 21.6 -2.785 21.7 -2.685 ;
        RECT 21.6 -3.775 21.7 -3.675 ;
        RECT 21.6 -4.13 21.7 -4.03 ;
        RECT 21.6 -5.66 21.7 -5.56 ;
        RECT 21.6 -6.015 21.7 -5.915 ;
        RECT 21.6 -7.005 21.7 -6.905 ;
        RECT 21.6 -7.36 21.7 -7.26 ;
        RECT 21.6 -8.89 21.7 -8.79 ;
        RECT 21.6 -9.245 21.7 -9.145 ;
        RECT 21.6 -10.235 21.7 -10.135 ;
        RECT 21.6 -10.59 21.7 -10.49 ;
        RECT 21.6 -12.12 21.7 -12.02 ;
        RECT 21.6 -12.475 21.7 -12.375 ;
        RECT 21.6 -13.465 21.7 -13.365 ;
        RECT 21.6 -13.82 21.7 -13.72 ;
        RECT 21.6 -15.35 21.7 -15.25 ;
        RECT 21.6 -15.705 21.7 -15.605 ;
        RECT 21.6 -16.695 21.7 -16.595 ;
        RECT 21.6 -17.05 21.7 -16.95 ;
        RECT 21.6 -18.58 21.7 -18.48 ;
        RECT 21.6 -18.935 21.7 -18.835 ;
        RECT 21.6 -19.925 21.7 -19.825 ;
        RECT 21.6 -20.28 21.7 -20.18 ;
        RECT 21.6 -21.81 21.7 -21.71 ;
        RECT 21.6 -22.165 21.7 -22.065 ;
        RECT 21.6 -23.155 21.7 -23.055 ;
        RECT 21.6 -23.51 21.7 -23.41 ;
        RECT 21.6 -25.04 21.7 -24.94 ;
        RECT 21.6 -25.395 21.7 -25.295 ;
        RECT 21.6 -26.385 21.7 -26.285 ;
        RECT 21.6 -26.74 21.7 -26.64 ;
        RECT 21.6 -28.27 21.7 -28.17 ;
        RECT 21.6 -28.625 21.7 -28.525 ;
        RECT 21.6 -29.615 21.7 -29.515 ;
        RECT 21.6 -29.97 21.7 -29.87 ;
        RECT 21.6 -31.5 21.7 -31.4 ;
        RECT 21.6 -31.855 21.7 -31.755 ;
        RECT 21.6 -32.845 21.7 -32.745 ;
        RECT 21.6 -33.2 21.7 -33.1 ;
        RECT 21.6 -34.73 21.7 -34.63 ;
        RECT 21.6 -35.085 21.7 -34.985 ;
        RECT 21.6 -36.075 21.7 -35.975 ;
        RECT 21.6 -36.43 21.7 -36.33 ;
        RECT 21.6 -37.96 21.7 -37.86 ;
        RECT 21.6 -38.315 21.7 -38.215 ;
        RECT 21.6 -39.305 21.7 -39.205 ;
        RECT 21.6 -39.66 21.7 -39.56 ;
        RECT 21.6 -41.19 21.7 -41.09 ;
        RECT 21.6 -41.545 21.7 -41.445 ;
        RECT 21.6 -42.535 21.7 -42.435 ;
        RECT 21.6 -42.89 21.7 -42.79 ;
        RECT 21.6 -44.42 21.7 -44.32 ;
        RECT 21.6 -44.775 21.7 -44.675 ;
        RECT 21.6 -45.765 21.7 -45.665 ;
        RECT 21.6 -46.12 21.7 -46.02 ;
        RECT 21.6 -47.65 21.7 -47.55 ;
        RECT 21.6 -48.005 21.7 -47.905 ;
        RECT 21.6 -48.995 21.7 -48.895 ;
        RECT 21.6 -49.35 21.7 -49.25 ;
        RECT 22.8 9.75 22.9 9.85 ;
        RECT 22.8 9.52 22.9 9.62 ;
        RECT 22.8 9.29 22.9 9.39 ;
        RECT 22.8 9.06 22.9 9.16 ;
        RECT 22.8 8.83 22.9 8.93 ;
        RECT 22.8 8.6 22.9 8.7 ;
        RECT 22.8 8.37 22.9 8.47 ;
        RECT 22.8 8.14 22.9 8.24 ;
        RECT 22.8 7.91 22.9 8.01 ;
        RECT 22.8 7.68 22.9 7.78 ;
        RECT 22.8 7.45 22.9 7.55 ;
        RECT 22.8 7.22 22.9 7.32 ;
        RECT 22.8 0.8 22.9 0.9 ;
        RECT 22.8 0.445 22.9 0.545 ;
        RECT 22.8 -0.545 22.9 -0.445 ;
        RECT 22.8 -0.9 22.9 -0.8 ;
        RECT 22.8 -2.43 22.9 -2.33 ;
        RECT 22.8 -2.785 22.9 -2.685 ;
        RECT 22.8 -3.775 22.9 -3.675 ;
        RECT 22.8 -4.13 22.9 -4.03 ;
        RECT 22.8 -5.66 22.9 -5.56 ;
        RECT 22.8 -6.015 22.9 -5.915 ;
        RECT 22.8 -7.005 22.9 -6.905 ;
        RECT 22.8 -7.36 22.9 -7.26 ;
        RECT 22.8 -8.89 22.9 -8.79 ;
        RECT 22.8 -9.245 22.9 -9.145 ;
        RECT 22.8 -10.235 22.9 -10.135 ;
        RECT 22.8 -10.59 22.9 -10.49 ;
        RECT 22.8 -12.12 22.9 -12.02 ;
        RECT 22.8 -12.475 22.9 -12.375 ;
        RECT 22.8 -13.465 22.9 -13.365 ;
        RECT 22.8 -13.82 22.9 -13.72 ;
        RECT 22.8 -15.35 22.9 -15.25 ;
        RECT 22.8 -15.705 22.9 -15.605 ;
        RECT 22.8 -16.695 22.9 -16.595 ;
        RECT 22.8 -17.05 22.9 -16.95 ;
        RECT 22.8 -18.58 22.9 -18.48 ;
        RECT 22.8 -18.935 22.9 -18.835 ;
        RECT 22.8 -19.925 22.9 -19.825 ;
        RECT 22.8 -20.28 22.9 -20.18 ;
        RECT 22.8 -21.81 22.9 -21.71 ;
        RECT 22.8 -22.165 22.9 -22.065 ;
        RECT 22.8 -23.155 22.9 -23.055 ;
        RECT 22.8 -23.51 22.9 -23.41 ;
        RECT 22.8 -25.04 22.9 -24.94 ;
        RECT 22.8 -25.395 22.9 -25.295 ;
        RECT 22.8 -26.385 22.9 -26.285 ;
        RECT 22.8 -26.74 22.9 -26.64 ;
        RECT 22.8 -28.27 22.9 -28.17 ;
        RECT 22.8 -28.625 22.9 -28.525 ;
        RECT 22.8 -29.615 22.9 -29.515 ;
        RECT 22.8 -29.97 22.9 -29.87 ;
        RECT 22.8 -31.5 22.9 -31.4 ;
        RECT 22.8 -31.855 22.9 -31.755 ;
        RECT 22.8 -32.845 22.9 -32.745 ;
        RECT 22.8 -33.2 22.9 -33.1 ;
        RECT 22.8 -34.73 22.9 -34.63 ;
        RECT 22.8 -35.085 22.9 -34.985 ;
        RECT 22.8 -36.075 22.9 -35.975 ;
        RECT 22.8 -36.43 22.9 -36.33 ;
        RECT 22.8 -37.96 22.9 -37.86 ;
        RECT 22.8 -38.315 22.9 -38.215 ;
        RECT 22.8 -39.305 22.9 -39.205 ;
        RECT 22.8 -39.66 22.9 -39.56 ;
        RECT 22.8 -41.19 22.9 -41.09 ;
        RECT 22.8 -41.545 22.9 -41.445 ;
        RECT 22.8 -42.535 22.9 -42.435 ;
        RECT 22.8 -42.89 22.9 -42.79 ;
        RECT 22.8 -44.42 22.9 -44.32 ;
        RECT 22.8 -44.775 22.9 -44.675 ;
        RECT 22.8 -45.765 22.9 -45.665 ;
        RECT 22.8 -46.12 22.9 -46.02 ;
        RECT 22.8 -47.65 22.9 -47.55 ;
        RECT 22.8 -48.005 22.9 -47.905 ;
        RECT 22.8 -48.995 22.9 -48.895 ;
        RECT 22.8 -49.35 22.9 -49.25 ;
        RECT 24 9.75 24.1 9.85 ;
        RECT 24 9.52 24.1 9.62 ;
        RECT 24 9.29 24.1 9.39 ;
        RECT 24 9.06 24.1 9.16 ;
        RECT 24 8.83 24.1 8.93 ;
        RECT 24 8.6 24.1 8.7 ;
        RECT 24 8.37 24.1 8.47 ;
        RECT 24 8.14 24.1 8.24 ;
        RECT 24 7.91 24.1 8.01 ;
        RECT 24 7.68 24.1 7.78 ;
        RECT 24 7.45 24.1 7.55 ;
        RECT 24 7.22 24.1 7.32 ;
        RECT 24 0.8 24.1 0.9 ;
        RECT 24 0.445 24.1 0.545 ;
        RECT 24 -0.545 24.1 -0.445 ;
        RECT 24 -0.9 24.1 -0.8 ;
        RECT 24 -2.43 24.1 -2.33 ;
        RECT 24 -2.785 24.1 -2.685 ;
        RECT 24 -3.775 24.1 -3.675 ;
        RECT 24 -4.13 24.1 -4.03 ;
        RECT 24 -5.66 24.1 -5.56 ;
        RECT 24 -6.015 24.1 -5.915 ;
        RECT 24 -7.005 24.1 -6.905 ;
        RECT 24 -7.36 24.1 -7.26 ;
        RECT 24 -8.89 24.1 -8.79 ;
        RECT 24 -9.245 24.1 -9.145 ;
        RECT 24 -10.235 24.1 -10.135 ;
        RECT 24 -10.59 24.1 -10.49 ;
        RECT 24 -12.12 24.1 -12.02 ;
        RECT 24 -12.475 24.1 -12.375 ;
        RECT 24 -13.465 24.1 -13.365 ;
        RECT 24 -13.82 24.1 -13.72 ;
        RECT 24 -15.35 24.1 -15.25 ;
        RECT 24 -15.705 24.1 -15.605 ;
        RECT 24 -16.695 24.1 -16.595 ;
        RECT 24 -17.05 24.1 -16.95 ;
        RECT 24 -18.58 24.1 -18.48 ;
        RECT 24 -18.935 24.1 -18.835 ;
        RECT 24 -19.925 24.1 -19.825 ;
        RECT 24 -20.28 24.1 -20.18 ;
        RECT 24 -21.81 24.1 -21.71 ;
        RECT 24 -22.165 24.1 -22.065 ;
        RECT 24 -23.155 24.1 -23.055 ;
        RECT 24 -23.51 24.1 -23.41 ;
        RECT 24 -25.04 24.1 -24.94 ;
        RECT 24 -25.395 24.1 -25.295 ;
        RECT 24 -26.385 24.1 -26.285 ;
        RECT 24 -26.74 24.1 -26.64 ;
        RECT 24 -28.27 24.1 -28.17 ;
        RECT 24 -28.625 24.1 -28.525 ;
        RECT 24 -29.615 24.1 -29.515 ;
        RECT 24 -29.97 24.1 -29.87 ;
        RECT 24 -31.5 24.1 -31.4 ;
        RECT 24 -31.855 24.1 -31.755 ;
        RECT 24 -32.845 24.1 -32.745 ;
        RECT 24 -33.2 24.1 -33.1 ;
        RECT 24 -34.73 24.1 -34.63 ;
        RECT 24 -35.085 24.1 -34.985 ;
        RECT 24 -36.075 24.1 -35.975 ;
        RECT 24 -36.43 24.1 -36.33 ;
        RECT 24 -37.96 24.1 -37.86 ;
        RECT 24 -38.315 24.1 -38.215 ;
        RECT 24 -39.305 24.1 -39.205 ;
        RECT 24 -39.66 24.1 -39.56 ;
        RECT 24 -41.19 24.1 -41.09 ;
        RECT 24 -41.545 24.1 -41.445 ;
        RECT 24 -42.535 24.1 -42.435 ;
        RECT 24 -42.89 24.1 -42.79 ;
        RECT 24 -44.42 24.1 -44.32 ;
        RECT 24 -44.775 24.1 -44.675 ;
        RECT 24 -45.765 24.1 -45.665 ;
        RECT 24 -46.12 24.1 -46.02 ;
        RECT 24 -47.65 24.1 -47.55 ;
        RECT 24 -48.005 24.1 -47.905 ;
        RECT 24 -48.995 24.1 -48.895 ;
        RECT 24 -49.35 24.1 -49.25 ;
        RECT 25.2 9.75 25.3 9.85 ;
        RECT 25.2 9.52 25.3 9.62 ;
        RECT 25.2 9.29 25.3 9.39 ;
        RECT 25.2 9.06 25.3 9.16 ;
        RECT 25.2 8.83 25.3 8.93 ;
        RECT 25.2 8.6 25.3 8.7 ;
        RECT 25.2 8.37 25.3 8.47 ;
        RECT 25.2 8.14 25.3 8.24 ;
        RECT 25.2 7.91 25.3 8.01 ;
        RECT 25.2 7.68 25.3 7.78 ;
        RECT 25.2 7.45 25.3 7.55 ;
        RECT 25.2 7.22 25.3 7.32 ;
        RECT 25.2 0.8 25.3 0.9 ;
        RECT 25.2 0.445 25.3 0.545 ;
        RECT 25.2 -0.545 25.3 -0.445 ;
        RECT 25.2 -0.9 25.3 -0.8 ;
        RECT 25.2 -2.43 25.3 -2.33 ;
        RECT 25.2 -2.785 25.3 -2.685 ;
        RECT 25.2 -3.775 25.3 -3.675 ;
        RECT 25.2 -4.13 25.3 -4.03 ;
        RECT 25.2 -5.66 25.3 -5.56 ;
        RECT 25.2 -6.015 25.3 -5.915 ;
        RECT 25.2 -7.005 25.3 -6.905 ;
        RECT 25.2 -7.36 25.3 -7.26 ;
        RECT 25.2 -8.89 25.3 -8.79 ;
        RECT 25.2 -9.245 25.3 -9.145 ;
        RECT 25.2 -10.235 25.3 -10.135 ;
        RECT 25.2 -10.59 25.3 -10.49 ;
        RECT 25.2 -12.12 25.3 -12.02 ;
        RECT 25.2 -12.475 25.3 -12.375 ;
        RECT 25.2 -13.465 25.3 -13.365 ;
        RECT 25.2 -13.82 25.3 -13.72 ;
        RECT 25.2 -15.35 25.3 -15.25 ;
        RECT 25.2 -15.705 25.3 -15.605 ;
        RECT 25.2 -16.695 25.3 -16.595 ;
        RECT 25.2 -17.05 25.3 -16.95 ;
        RECT 25.2 -18.58 25.3 -18.48 ;
        RECT 25.2 -18.935 25.3 -18.835 ;
        RECT 25.2 -19.925 25.3 -19.825 ;
        RECT 25.2 -20.28 25.3 -20.18 ;
        RECT 25.2 -21.81 25.3 -21.71 ;
        RECT 25.2 -22.165 25.3 -22.065 ;
        RECT 25.2 -23.155 25.3 -23.055 ;
        RECT 25.2 -23.51 25.3 -23.41 ;
        RECT 25.2 -25.04 25.3 -24.94 ;
        RECT 25.2 -25.395 25.3 -25.295 ;
        RECT 25.2 -26.385 25.3 -26.285 ;
        RECT 25.2 -26.74 25.3 -26.64 ;
        RECT 25.2 -28.27 25.3 -28.17 ;
        RECT 25.2 -28.625 25.3 -28.525 ;
        RECT 25.2 -29.615 25.3 -29.515 ;
        RECT 25.2 -29.97 25.3 -29.87 ;
        RECT 25.2 -31.5 25.3 -31.4 ;
        RECT 25.2 -31.855 25.3 -31.755 ;
        RECT 25.2 -32.845 25.3 -32.745 ;
        RECT 25.2 -33.2 25.3 -33.1 ;
        RECT 25.2 -34.73 25.3 -34.63 ;
        RECT 25.2 -35.085 25.3 -34.985 ;
        RECT 25.2 -36.075 25.3 -35.975 ;
        RECT 25.2 -36.43 25.3 -36.33 ;
        RECT 25.2 -37.96 25.3 -37.86 ;
        RECT 25.2 -38.315 25.3 -38.215 ;
        RECT 25.2 -39.305 25.3 -39.205 ;
        RECT 25.2 -39.66 25.3 -39.56 ;
        RECT 25.2 -41.19 25.3 -41.09 ;
        RECT 25.2 -41.545 25.3 -41.445 ;
        RECT 25.2 -42.535 25.3 -42.435 ;
        RECT 25.2 -42.89 25.3 -42.79 ;
        RECT 25.2 -44.42 25.3 -44.32 ;
        RECT 25.2 -44.775 25.3 -44.675 ;
        RECT 25.2 -45.765 25.3 -45.665 ;
        RECT 25.2 -46.12 25.3 -46.02 ;
        RECT 25.2 -47.65 25.3 -47.55 ;
        RECT 25.2 -48.005 25.3 -47.905 ;
        RECT 25.2 -48.995 25.3 -48.895 ;
        RECT 25.2 -49.35 25.3 -49.25 ;
        RECT 26.4 9.75 26.5 9.85 ;
        RECT 26.4 9.52 26.5 9.62 ;
        RECT 26.4 9.29 26.5 9.39 ;
        RECT 26.4 9.06 26.5 9.16 ;
        RECT 26.4 8.83 26.5 8.93 ;
        RECT 26.4 8.6 26.5 8.7 ;
        RECT 26.4 8.37 26.5 8.47 ;
        RECT 26.4 8.14 26.5 8.24 ;
        RECT 26.4 7.91 26.5 8.01 ;
        RECT 26.4 7.68 26.5 7.78 ;
        RECT 26.4 7.45 26.5 7.55 ;
        RECT 26.4 7.22 26.5 7.32 ;
        RECT 26.4 0.8 26.5 0.9 ;
        RECT 26.4 0.445 26.5 0.545 ;
        RECT 26.4 -0.545 26.5 -0.445 ;
        RECT 26.4 -0.9 26.5 -0.8 ;
        RECT 26.4 -2.43 26.5 -2.33 ;
        RECT 26.4 -2.785 26.5 -2.685 ;
        RECT 26.4 -3.775 26.5 -3.675 ;
        RECT 26.4 -4.13 26.5 -4.03 ;
        RECT 26.4 -5.66 26.5 -5.56 ;
        RECT 26.4 -6.015 26.5 -5.915 ;
        RECT 26.4 -7.005 26.5 -6.905 ;
        RECT 26.4 -7.36 26.5 -7.26 ;
        RECT 26.4 -8.89 26.5 -8.79 ;
        RECT 26.4 -9.245 26.5 -9.145 ;
        RECT 26.4 -10.235 26.5 -10.135 ;
        RECT 26.4 -10.59 26.5 -10.49 ;
        RECT 26.4 -12.12 26.5 -12.02 ;
        RECT 26.4 -12.475 26.5 -12.375 ;
        RECT 26.4 -13.465 26.5 -13.365 ;
        RECT 26.4 -13.82 26.5 -13.72 ;
        RECT 26.4 -15.35 26.5 -15.25 ;
        RECT 26.4 -15.705 26.5 -15.605 ;
        RECT 26.4 -16.695 26.5 -16.595 ;
        RECT 26.4 -17.05 26.5 -16.95 ;
        RECT 26.4 -18.58 26.5 -18.48 ;
        RECT 26.4 -18.935 26.5 -18.835 ;
        RECT 26.4 -19.925 26.5 -19.825 ;
        RECT 26.4 -20.28 26.5 -20.18 ;
        RECT 26.4 -21.81 26.5 -21.71 ;
        RECT 26.4 -22.165 26.5 -22.065 ;
        RECT 26.4 -23.155 26.5 -23.055 ;
        RECT 26.4 -23.51 26.5 -23.41 ;
        RECT 26.4 -25.04 26.5 -24.94 ;
        RECT 26.4 -25.395 26.5 -25.295 ;
        RECT 26.4 -26.385 26.5 -26.285 ;
        RECT 26.4 -26.74 26.5 -26.64 ;
        RECT 26.4 -28.27 26.5 -28.17 ;
        RECT 26.4 -28.625 26.5 -28.525 ;
        RECT 26.4 -29.615 26.5 -29.515 ;
        RECT 26.4 -29.97 26.5 -29.87 ;
        RECT 26.4 -31.5 26.5 -31.4 ;
        RECT 26.4 -31.855 26.5 -31.755 ;
        RECT 26.4 -32.845 26.5 -32.745 ;
        RECT 26.4 -33.2 26.5 -33.1 ;
        RECT 26.4 -34.73 26.5 -34.63 ;
        RECT 26.4 -35.085 26.5 -34.985 ;
        RECT 26.4 -36.075 26.5 -35.975 ;
        RECT 26.4 -36.43 26.5 -36.33 ;
        RECT 26.4 -37.96 26.5 -37.86 ;
        RECT 26.4 -38.315 26.5 -38.215 ;
        RECT 26.4 -39.305 26.5 -39.205 ;
        RECT 26.4 -39.66 26.5 -39.56 ;
        RECT 26.4 -41.19 26.5 -41.09 ;
        RECT 26.4 -41.545 26.5 -41.445 ;
        RECT 26.4 -42.535 26.5 -42.435 ;
        RECT 26.4 -42.89 26.5 -42.79 ;
        RECT 26.4 -44.42 26.5 -44.32 ;
        RECT 26.4 -44.775 26.5 -44.675 ;
        RECT 26.4 -45.765 26.5 -45.665 ;
        RECT 26.4 -46.12 26.5 -46.02 ;
        RECT 26.4 -47.65 26.5 -47.55 ;
        RECT 26.4 -48.005 26.5 -47.905 ;
        RECT 26.4 -48.995 26.5 -48.895 ;
        RECT 26.4 -49.35 26.5 -49.25 ;
        RECT 27.6 9.75 27.7 9.85 ;
        RECT 27.6 9.52 27.7 9.62 ;
        RECT 27.6 9.29 27.7 9.39 ;
        RECT 27.6 9.06 27.7 9.16 ;
        RECT 27.6 8.83 27.7 8.93 ;
        RECT 27.6 8.6 27.7 8.7 ;
        RECT 27.6 8.37 27.7 8.47 ;
        RECT 27.6 8.14 27.7 8.24 ;
        RECT 27.6 7.91 27.7 8.01 ;
        RECT 27.6 7.68 27.7 7.78 ;
        RECT 27.6 7.45 27.7 7.55 ;
        RECT 27.6 7.22 27.7 7.32 ;
        RECT 27.6 0.8 27.7 0.9 ;
        RECT 27.6 0.445 27.7 0.545 ;
        RECT 27.6 -0.545 27.7 -0.445 ;
        RECT 27.6 -0.9 27.7 -0.8 ;
        RECT 27.6 -2.43 27.7 -2.33 ;
        RECT 27.6 -2.785 27.7 -2.685 ;
        RECT 27.6 -3.775 27.7 -3.675 ;
        RECT 27.6 -4.13 27.7 -4.03 ;
        RECT 27.6 -5.66 27.7 -5.56 ;
        RECT 27.6 -6.015 27.7 -5.915 ;
        RECT 27.6 -7.005 27.7 -6.905 ;
        RECT 27.6 -7.36 27.7 -7.26 ;
        RECT 27.6 -8.89 27.7 -8.79 ;
        RECT 27.6 -9.245 27.7 -9.145 ;
        RECT 27.6 -10.235 27.7 -10.135 ;
        RECT 27.6 -10.59 27.7 -10.49 ;
        RECT 27.6 -12.12 27.7 -12.02 ;
        RECT 27.6 -12.475 27.7 -12.375 ;
        RECT 27.6 -13.465 27.7 -13.365 ;
        RECT 27.6 -13.82 27.7 -13.72 ;
        RECT 27.6 -15.35 27.7 -15.25 ;
        RECT 27.6 -15.705 27.7 -15.605 ;
        RECT 27.6 -16.695 27.7 -16.595 ;
        RECT 27.6 -17.05 27.7 -16.95 ;
        RECT 27.6 -18.58 27.7 -18.48 ;
        RECT 27.6 -18.935 27.7 -18.835 ;
        RECT 27.6 -19.925 27.7 -19.825 ;
        RECT 27.6 -20.28 27.7 -20.18 ;
        RECT 27.6 -21.81 27.7 -21.71 ;
        RECT 27.6 -22.165 27.7 -22.065 ;
        RECT 27.6 -23.155 27.7 -23.055 ;
        RECT 27.6 -23.51 27.7 -23.41 ;
        RECT 27.6 -25.04 27.7 -24.94 ;
        RECT 27.6 -25.395 27.7 -25.295 ;
        RECT 27.6 -26.385 27.7 -26.285 ;
        RECT 27.6 -26.74 27.7 -26.64 ;
        RECT 27.6 -28.27 27.7 -28.17 ;
        RECT 27.6 -28.625 27.7 -28.525 ;
        RECT 27.6 -29.615 27.7 -29.515 ;
        RECT 27.6 -29.97 27.7 -29.87 ;
        RECT 27.6 -31.5 27.7 -31.4 ;
        RECT 27.6 -31.855 27.7 -31.755 ;
        RECT 27.6 -32.845 27.7 -32.745 ;
        RECT 27.6 -33.2 27.7 -33.1 ;
        RECT 27.6 -34.73 27.7 -34.63 ;
        RECT 27.6 -35.085 27.7 -34.985 ;
        RECT 27.6 -36.075 27.7 -35.975 ;
        RECT 27.6 -36.43 27.7 -36.33 ;
        RECT -33.42 9.75 -33.32 9.85 ;
        RECT -33.42 9.52 -33.32 9.62 ;
        RECT -33.42 9.29 -33.32 9.39 ;
        RECT -33.42 9.06 -33.32 9.16 ;
        RECT -33.42 8.83 -33.32 8.93 ;
        RECT -33.42 8.6 -33.32 8.7 ;
        RECT -33.42 8.37 -33.32 8.47 ;
        RECT -33.42 8.14 -33.32 8.24 ;
        RECT -33.42 7.91 -33.32 8.01 ;
        RECT -33.42 7.68 -33.32 7.78 ;
        RECT -33.42 7.45 -33.32 7.55 ;
        RECT -33.42 7.22 -33.32 7.32 ;
        RECT -33.42 5.795 -33.32 5.895 ;
        RECT -33.42 5.565 -33.32 5.665 ;
        RECT -33.42 5.335 -33.32 5.435 ;
        RECT -33.42 -4.665 -33.32 -4.565 ;
        RECT -33.42 -4.895 -33.32 -4.795 ;
        RECT -33.42 -5.125 -33.32 -5.025 ;
        RECT -33.42 -17.585 -33.32 -17.485 ;
        RECT -33.42 -17.815 -33.32 -17.715 ;
        RECT -33.42 -18.045 -33.32 -17.945 ;
        RECT -33.42 -30.505 -33.32 -30.405 ;
        RECT -33.42 -30.735 -33.32 -30.635 ;
        RECT -33.42 -30.965 -33.32 -30.865 ;
        RECT -33.42 -43.425 -33.32 -43.325 ;
        RECT -33.42 -43.655 -33.32 -43.555 ;
        RECT -33.42 -43.885 -33.32 -43.785 ;
        RECT -33.42 -56.345 -33.32 -56.245 ;
        RECT -33.42 -56.575 -33.32 -56.475 ;
        RECT -33.42 -56.805 -33.32 -56.705 ;
        RECT -33.19 9.75 -33.09 9.85 ;
        RECT -33.19 9.52 -33.09 9.62 ;
        RECT -33.19 9.29 -33.09 9.39 ;
        RECT -33.19 9.06 -33.09 9.16 ;
        RECT -33.19 8.83 -33.09 8.93 ;
        RECT -33.19 8.6 -33.09 8.7 ;
        RECT -33.19 8.37 -33.09 8.47 ;
        RECT -33.19 8.14 -33.09 8.24 ;
        RECT -33.19 7.91 -33.09 8.01 ;
        RECT -33.19 7.68 -33.09 7.78 ;
        RECT -33.19 7.45 -33.09 7.55 ;
        RECT -33.19 7.22 -33.09 7.32 ;
        RECT -33.19 5.795 -33.09 5.895 ;
        RECT -33.19 5.565 -33.09 5.665 ;
        RECT -33.19 5.335 -33.09 5.435 ;
        RECT -33.19 -4.665 -33.09 -4.565 ;
        RECT -33.19 -4.895 -33.09 -4.795 ;
        RECT -33.19 -5.125 -33.09 -5.025 ;
        RECT -33.19 -17.585 -33.09 -17.485 ;
        RECT -33.19 -17.815 -33.09 -17.715 ;
        RECT -33.19 -18.045 -33.09 -17.945 ;
        RECT -33.19 -30.505 -33.09 -30.405 ;
        RECT -33.19 -30.735 -33.09 -30.635 ;
        RECT -33.19 -30.965 -33.09 -30.865 ;
        RECT -33.19 -43.425 -33.09 -43.325 ;
        RECT -33.19 -43.655 -33.09 -43.555 ;
        RECT -33.19 -43.885 -33.09 -43.785 ;
        RECT -33.19 -56.345 -33.09 -56.245 ;
        RECT -33.19 -56.575 -33.09 -56.475 ;
        RECT -33.19 -56.805 -33.09 -56.705 ;
        RECT -32.96 9.75 -32.86 9.85 ;
        RECT -32.96 9.52 -32.86 9.62 ;
        RECT -32.96 9.29 -32.86 9.39 ;
        RECT -32.96 9.06 -32.86 9.16 ;
        RECT -32.96 8.83 -32.86 8.93 ;
        RECT -32.96 8.6 -32.86 8.7 ;
        RECT -32.96 8.37 -32.86 8.47 ;
        RECT -32.96 8.14 -32.86 8.24 ;
        RECT -32.96 7.91 -32.86 8.01 ;
        RECT -32.96 7.68 -32.86 7.78 ;
        RECT -32.96 7.45 -32.86 7.55 ;
        RECT -32.96 7.22 -32.86 7.32 ;
        RECT -32.96 5.795 -32.86 5.895 ;
        RECT -32.96 5.565 -32.86 5.665 ;
        RECT -32.96 5.335 -32.86 5.435 ;
        RECT -32.96 -4.665 -32.86 -4.565 ;
        RECT -32.96 -4.895 -32.86 -4.795 ;
        RECT -32.96 -5.125 -32.86 -5.025 ;
        RECT -32.96 -17.585 -32.86 -17.485 ;
        RECT -32.96 -17.815 -32.86 -17.715 ;
        RECT -32.96 -18.045 -32.86 -17.945 ;
        RECT -32.96 -30.505 -32.86 -30.405 ;
        RECT -32.96 -30.735 -32.86 -30.635 ;
        RECT -32.96 -30.965 -32.86 -30.865 ;
        RECT -32.96 -43.425 -32.86 -43.325 ;
        RECT -32.96 -43.655 -32.86 -43.555 ;
        RECT -32.96 -43.885 -32.86 -43.785 ;
        RECT -32.96 -56.345 -32.86 -56.245 ;
        RECT -32.96 -56.575 -32.86 -56.475 ;
        RECT -32.96 -56.805 -32.86 -56.705 ;
        RECT -32.73 9.75 -32.63 9.85 ;
        RECT -32.73 9.52 -32.63 9.62 ;
        RECT -32.73 9.29 -32.63 9.39 ;
        RECT -32.73 9.06 -32.63 9.16 ;
        RECT -32.73 8.83 -32.63 8.93 ;
        RECT -32.73 8.6 -32.63 8.7 ;
        RECT -32.73 8.37 -32.63 8.47 ;
        RECT -32.73 8.14 -32.63 8.24 ;
        RECT -32.73 7.91 -32.63 8.01 ;
        RECT -32.73 7.68 -32.63 7.78 ;
        RECT -32.73 7.45 -32.63 7.55 ;
        RECT -32.73 7.22 -32.63 7.32 ;
        RECT -32.73 5.795 -32.63 5.895 ;
        RECT -32.73 5.565 -32.63 5.665 ;
        RECT -32.73 5.335 -32.63 5.435 ;
        RECT -32.73 -4.665 -32.63 -4.565 ;
        RECT -32.73 -4.895 -32.63 -4.795 ;
        RECT -32.73 -5.125 -32.63 -5.025 ;
        RECT -32.73 -17.585 -32.63 -17.485 ;
        RECT -32.73 -17.815 -32.63 -17.715 ;
        RECT -32.73 -18.045 -32.63 -17.945 ;
        RECT -32.73 -30.505 -32.63 -30.405 ;
        RECT -32.73 -30.735 -32.63 -30.635 ;
        RECT -32.73 -30.965 -32.63 -30.865 ;
        RECT -32.73 -43.425 -32.63 -43.325 ;
        RECT -32.73 -43.655 -32.63 -43.555 ;
        RECT -32.73 -43.885 -32.63 -43.785 ;
        RECT -32.73 -56.345 -32.63 -56.245 ;
        RECT -32.73 -56.575 -32.63 -56.475 ;
        RECT -32.73 -56.805 -32.63 -56.705 ;
        RECT -5.705 -3.985 -5.605 -3.885 ;
        RECT -5.705 -4.225 -5.605 -4.125 ;
        RECT -5.705 -5.565 -5.605 -5.465 ;
        RECT -5.705 -5.805 -5.605 -5.705 ;
        RECT -5.705 -16.905 -5.605 -16.805 ;
        RECT -5.705 -17.145 -5.605 -17.045 ;
        RECT -5.705 -18.485 -5.605 -18.385 ;
        RECT -5.705 -18.725 -5.605 -18.625 ;
        RECT -5.705 -29.825 -5.605 -29.725 ;
        RECT -5.705 -30.065 -5.605 -29.965 ;
        RECT -5.705 -31.405 -5.605 -31.305 ;
        RECT -5.705 -31.645 -5.605 -31.545 ;
        RECT -5.705 -42.745 -5.605 -42.645 ;
        RECT -5.705 -42.985 -5.605 -42.885 ;
        RECT -5.705 -44.325 -5.605 -44.225 ;
        RECT -5.705 -44.565 -5.605 -44.465 ;
        RECT -5.705 -55.665 -5.605 -55.565 ;
        RECT -5.705 -55.905 -5.605 -55.805 ;
        RECT -4.405 -3.985 -4.305 -3.885 ;
        RECT -4.405 -4.225 -4.305 -4.125 ;
        RECT -4.405 -5.565 -4.305 -5.465 ;
        RECT -4.405 -5.805 -4.305 -5.705 ;
        RECT -4.405 -16.905 -4.305 -16.805 ;
        RECT -4.405 -17.145 -4.305 -17.045 ;
        RECT -4.405 -18.485 -4.305 -18.385 ;
        RECT -4.405 -18.725 -4.305 -18.625 ;
        RECT -4.405 -29.825 -4.305 -29.725 ;
        RECT -4.405 -30.065 -4.305 -29.965 ;
        RECT -4.405 -31.405 -4.305 -31.305 ;
        RECT -4.405 -31.645 -4.305 -31.545 ;
        RECT -4.405 -42.745 -4.305 -42.645 ;
        RECT -4.405 -42.985 -4.305 -42.885 ;
        RECT -4.405 -44.325 -4.305 -44.225 ;
        RECT -4.405 -44.565 -4.305 -44.465 ;
        RECT -4.405 -55.665 -4.305 -55.565 ;
        RECT -4.405 -55.905 -4.305 -55.805 ;
        RECT -3.105 -3.985 -3.005 -3.885 ;
        RECT -3.105 -4.225 -3.005 -4.125 ;
        RECT -3.105 -5.565 -3.005 -5.465 ;
        RECT -3.105 -5.805 -3.005 -5.705 ;
        RECT -3.105 -16.905 -3.005 -16.805 ;
        RECT -3.105 -17.145 -3.005 -17.045 ;
        RECT -3.105 -18.485 -3.005 -18.385 ;
        RECT -3.105 -18.725 -3.005 -18.625 ;
        RECT -3.105 -29.825 -3.005 -29.725 ;
        RECT -3.105 -30.065 -3.005 -29.965 ;
        RECT -3.105 -31.405 -3.005 -31.305 ;
        RECT -3.105 -31.645 -3.005 -31.545 ;
        RECT -3.105 -42.745 -3.005 -42.645 ;
        RECT -3.105 -42.985 -3.005 -42.885 ;
        RECT -3.105 -44.325 -3.005 -44.225 ;
        RECT -3.105 -44.565 -3.005 -44.465 ;
        RECT -3.105 -55.665 -3.005 -55.565 ;
        RECT -3.105 -55.905 -3.005 -55.805 ;
        RECT -1.805 -3.985 -1.705 -3.885 ;
        RECT -1.805 -4.225 -1.705 -4.125 ;
        RECT -1.805 -5.565 -1.705 -5.465 ;
        RECT -1.805 -5.805 -1.705 -5.705 ;
        RECT -1.805 -16.905 -1.705 -16.805 ;
        RECT -1.805 -17.145 -1.705 -17.045 ;
        RECT -1.805 -18.485 -1.705 -18.385 ;
        RECT -1.805 -18.725 -1.705 -18.625 ;
        RECT -1.805 -29.825 -1.705 -29.725 ;
        RECT -1.805 -30.065 -1.705 -29.965 ;
        RECT -1.805 -31.405 -1.705 -31.305 ;
        RECT -1.805 -31.645 -1.705 -31.545 ;
        RECT -1.805 -42.745 -1.705 -42.645 ;
        RECT -1.805 -42.985 -1.705 -42.885 ;
        RECT -1.805 -44.325 -1.705 -44.225 ;
        RECT -1.805 -44.565 -1.705 -44.465 ;
        RECT -1.805 -55.665 -1.705 -55.565 ;
        RECT -1.805 -55.905 -1.705 -55.805 ;
        RECT 0 9.75 0.1 9.85 ;
        RECT 0 9.52 0.1 9.62 ;
        RECT 0 9.29 0.1 9.39 ;
        RECT 0 9.06 0.1 9.16 ;
        RECT 0 8.83 0.1 8.93 ;
        RECT 0 8.6 0.1 8.7 ;
        RECT 0 8.37 0.1 8.47 ;
        RECT 0 8.14 0.1 8.24 ;
        RECT 0 7.91 0.1 8.01 ;
        RECT 0 7.68 0.1 7.78 ;
        RECT 0 7.45 0.1 7.55 ;
        RECT 0 7.22 0.1 7.32 ;
        RECT 0 0.8 0.1 0.9 ;
        RECT 0 0.445 0.1 0.545 ;
        RECT 0 -0.545 0.1 -0.445 ;
        RECT 0 -0.9 0.1 -0.8 ;
        RECT 0 -2.43 0.1 -2.33 ;
        RECT 0 -2.785 0.1 -2.685 ;
        RECT 0 -3.775 0.1 -3.675 ;
        RECT 0 -4.13 0.1 -4.03 ;
        RECT 0 -5.66 0.1 -5.56 ;
        RECT 0 -6.015 0.1 -5.915 ;
        RECT 0 -7.005 0.1 -6.905 ;
        RECT 0 -7.36 0.1 -7.26 ;
        RECT 0 -8.89 0.1 -8.79 ;
        RECT 0 -9.245 0.1 -9.145 ;
        RECT 0 -10.235 0.1 -10.135 ;
        RECT 0 -10.59 0.1 -10.49 ;
        RECT 0 -12.12 0.1 -12.02 ;
        RECT 0 -12.475 0.1 -12.375 ;
        RECT 0 -13.465 0.1 -13.365 ;
        RECT 0 -13.82 0.1 -13.72 ;
        RECT 0 -15.35 0.1 -15.25 ;
        RECT 0 -15.705 0.1 -15.605 ;
        RECT 0 -16.695 0.1 -16.595 ;
        RECT 0 -17.05 0.1 -16.95 ;
        RECT 0 -18.58 0.1 -18.48 ;
        RECT 0 -18.935 0.1 -18.835 ;
        RECT 0 -19.925 0.1 -19.825 ;
        RECT 0 -20.28 0.1 -20.18 ;
        RECT 0 -21.81 0.1 -21.71 ;
        RECT 0 -22.165 0.1 -22.065 ;
        RECT 0 -23.155 0.1 -23.055 ;
        RECT 0 -23.51 0.1 -23.41 ;
        RECT 0 -25.04 0.1 -24.94 ;
        RECT 0 -25.395 0.1 -25.295 ;
        RECT 0 -26.385 0.1 -26.285 ;
        RECT 0 -26.74 0.1 -26.64 ;
        RECT 0 -28.27 0.1 -28.17 ;
        RECT 0 -28.625 0.1 -28.525 ;
        RECT 0 -29.615 0.1 -29.515 ;
        RECT 0 -29.97 0.1 -29.87 ;
        RECT 0 -31.5 0.1 -31.4 ;
        RECT 0 -31.855 0.1 -31.755 ;
        RECT 0 -32.845 0.1 -32.745 ;
        RECT 0 -33.2 0.1 -33.1 ;
        RECT 0 -34.73 0.1 -34.63 ;
        RECT 0 -35.085 0.1 -34.985 ;
        RECT 0 -36.075 0.1 -35.975 ;
        RECT 0 -36.43 0.1 -36.33 ;
        RECT 0 -37.96 0.1 -37.86 ;
        RECT 0 -38.315 0.1 -38.215 ;
        RECT 0 -39.305 0.1 -39.205 ;
        RECT 0 -39.66 0.1 -39.56 ;
        RECT 0 -41.19 0.1 -41.09 ;
        RECT 0 -41.545 0.1 -41.445 ;
        RECT 0 -42.535 0.1 -42.435 ;
        RECT 0 -42.89 0.1 -42.79 ;
        RECT 0 -44.42 0.1 -44.32 ;
        RECT 0 -44.775 0.1 -44.675 ;
        RECT 0 -45.765 0.1 -45.665 ;
        RECT 0 -46.12 0.1 -46.02 ;
        RECT 0 -47.65 0.1 -47.55 ;
        RECT 0 -48.005 0.1 -47.905 ;
        RECT 0 -48.995 0.1 -48.895 ;
        RECT 0 -49.35 0.1 -49.25 ;
        RECT 1.2 9.75 1.3 9.85 ;
        RECT 1.2 9.52 1.3 9.62 ;
        RECT 1.2 9.29 1.3 9.39 ;
        RECT 1.2 9.06 1.3 9.16 ;
        RECT 1.2 8.83 1.3 8.93 ;
        RECT 1.2 8.6 1.3 8.7 ;
        RECT 1.2 8.37 1.3 8.47 ;
        RECT 1.2 8.14 1.3 8.24 ;
        RECT 1.2 7.91 1.3 8.01 ;
        RECT 1.2 7.68 1.3 7.78 ;
        RECT 1.2 7.45 1.3 7.55 ;
        RECT 1.2 7.22 1.3 7.32 ;
        RECT 1.2 0.8 1.3 0.9 ;
        RECT 1.2 0.445 1.3 0.545 ;
        RECT 1.2 -0.545 1.3 -0.445 ;
        RECT 1.2 -0.9 1.3 -0.8 ;
        RECT 1.2 -2.43 1.3 -2.33 ;
        RECT 1.2 -2.785 1.3 -2.685 ;
        RECT 1.2 -3.775 1.3 -3.675 ;
        RECT 1.2 -4.13 1.3 -4.03 ;
        RECT 1.2 -5.66 1.3 -5.56 ;
        RECT 1.2 -6.015 1.3 -5.915 ;
        RECT 1.2 -7.005 1.3 -6.905 ;
        RECT 1.2 -7.36 1.3 -7.26 ;
        RECT 1.2 -8.89 1.3 -8.79 ;
        RECT 1.2 -9.245 1.3 -9.145 ;
        RECT 1.2 -10.235 1.3 -10.135 ;
        RECT 1.2 -10.59 1.3 -10.49 ;
        RECT 1.2 -12.12 1.3 -12.02 ;
        RECT 1.2 -12.475 1.3 -12.375 ;
        RECT 1.2 -13.465 1.3 -13.365 ;
        RECT 1.2 -13.82 1.3 -13.72 ;
        RECT 1.2 -15.35 1.3 -15.25 ;
        RECT 1.2 -15.705 1.3 -15.605 ;
        RECT 1.2 -16.695 1.3 -16.595 ;
        RECT 1.2 -17.05 1.3 -16.95 ;
        RECT 1.2 -18.58 1.3 -18.48 ;
        RECT 1.2 -18.935 1.3 -18.835 ;
        RECT 1.2 -19.925 1.3 -19.825 ;
        RECT 1.2 -20.28 1.3 -20.18 ;
        RECT 1.2 -21.81 1.3 -21.71 ;
        RECT 1.2 -22.165 1.3 -22.065 ;
        RECT 1.2 -23.155 1.3 -23.055 ;
        RECT 1.2 -23.51 1.3 -23.41 ;
        RECT 1.2 -25.04 1.3 -24.94 ;
        RECT 1.2 -25.395 1.3 -25.295 ;
        RECT 1.2 -26.385 1.3 -26.285 ;
        RECT 1.2 -26.74 1.3 -26.64 ;
        RECT 1.2 -28.27 1.3 -28.17 ;
        RECT 1.2 -28.625 1.3 -28.525 ;
        RECT 1.2 -29.615 1.3 -29.515 ;
        RECT 1.2 -29.97 1.3 -29.87 ;
        RECT 1.2 -31.5 1.3 -31.4 ;
        RECT 1.2 -31.855 1.3 -31.755 ;
        RECT 1.2 -32.845 1.3 -32.745 ;
        RECT 1.2 -33.2 1.3 -33.1 ;
        RECT 1.2 -34.73 1.3 -34.63 ;
        RECT 1.2 -35.085 1.3 -34.985 ;
        RECT 1.2 -36.075 1.3 -35.975 ;
        RECT 1.2 -36.43 1.3 -36.33 ;
        RECT 1.2 -37.96 1.3 -37.86 ;
        RECT 1.2 -38.315 1.3 -38.215 ;
        RECT 1.2 -39.305 1.3 -39.205 ;
        RECT 1.2 -39.66 1.3 -39.56 ;
        RECT 1.2 -41.19 1.3 -41.09 ;
        RECT 1.2 -41.545 1.3 -41.445 ;
        RECT 1.2 -42.535 1.3 -42.435 ;
        RECT 1.2 -42.89 1.3 -42.79 ;
        RECT 1.2 -44.42 1.3 -44.32 ;
        RECT 1.2 -44.775 1.3 -44.675 ;
        RECT 1.2 -45.765 1.3 -45.665 ;
        RECT 1.2 -46.12 1.3 -46.02 ;
        RECT 1.2 -47.65 1.3 -47.55 ;
        RECT 1.2 -48.005 1.3 -47.905 ;
        RECT 1.2 -48.995 1.3 -48.895 ;
        RECT 1.2 -49.35 1.3 -49.25 ;
        RECT 2.4 9.75 2.5 9.85 ;
        RECT 2.4 9.52 2.5 9.62 ;
        RECT 2.4 9.29 2.5 9.39 ;
        RECT 2.4 9.06 2.5 9.16 ;
        RECT 2.4 8.83 2.5 8.93 ;
        RECT 2.4 8.6 2.5 8.7 ;
        RECT 2.4 8.37 2.5 8.47 ;
        RECT 2.4 8.14 2.5 8.24 ;
        RECT 2.4 7.91 2.5 8.01 ;
        RECT 2.4 7.68 2.5 7.78 ;
        RECT 2.4 7.45 2.5 7.55 ;
        RECT 2.4 7.22 2.5 7.32 ;
        RECT 2.4 0.8 2.5 0.9 ;
        RECT 2.4 0.445 2.5 0.545 ;
        RECT 2.4 -0.545 2.5 -0.445 ;
        RECT 2.4 -0.9 2.5 -0.8 ;
        RECT 2.4 -2.43 2.5 -2.33 ;
        RECT 2.4 -2.785 2.5 -2.685 ;
        RECT 2.4 -3.775 2.5 -3.675 ;
        RECT 2.4 -4.13 2.5 -4.03 ;
        RECT 2.4 -5.66 2.5 -5.56 ;
        RECT 2.4 -6.015 2.5 -5.915 ;
        RECT 2.4 -7.005 2.5 -6.905 ;
        RECT 2.4 -7.36 2.5 -7.26 ;
        RECT 2.4 -8.89 2.5 -8.79 ;
        RECT 2.4 -9.245 2.5 -9.145 ;
        RECT 2.4 -10.235 2.5 -10.135 ;
        RECT 2.4 -10.59 2.5 -10.49 ;
        RECT 2.4 -12.12 2.5 -12.02 ;
        RECT 2.4 -12.475 2.5 -12.375 ;
        RECT 2.4 -13.465 2.5 -13.365 ;
        RECT 2.4 -13.82 2.5 -13.72 ;
        RECT 2.4 -15.35 2.5 -15.25 ;
        RECT 2.4 -15.705 2.5 -15.605 ;
        RECT 2.4 -16.695 2.5 -16.595 ;
        RECT 2.4 -17.05 2.5 -16.95 ;
        RECT 2.4 -18.58 2.5 -18.48 ;
        RECT 2.4 -18.935 2.5 -18.835 ;
        RECT 2.4 -19.925 2.5 -19.825 ;
        RECT 2.4 -20.28 2.5 -20.18 ;
        RECT 2.4 -21.81 2.5 -21.71 ;
        RECT 2.4 -22.165 2.5 -22.065 ;
        RECT 2.4 -23.155 2.5 -23.055 ;
        RECT 2.4 -23.51 2.5 -23.41 ;
        RECT 2.4 -25.04 2.5 -24.94 ;
        RECT 2.4 -25.395 2.5 -25.295 ;
        RECT 2.4 -26.385 2.5 -26.285 ;
        RECT 2.4 -26.74 2.5 -26.64 ;
        RECT 2.4 -28.27 2.5 -28.17 ;
        RECT 2.4 -28.625 2.5 -28.525 ;
        RECT 2.4 -29.615 2.5 -29.515 ;
        RECT 2.4 -29.97 2.5 -29.87 ;
        RECT 2.4 -31.5 2.5 -31.4 ;
        RECT 2.4 -31.855 2.5 -31.755 ;
        RECT 2.4 -32.845 2.5 -32.745 ;
        RECT 2.4 -33.2 2.5 -33.1 ;
        RECT 2.4 -34.73 2.5 -34.63 ;
        RECT 2.4 -35.085 2.5 -34.985 ;
        RECT 2.4 -36.075 2.5 -35.975 ;
        RECT 2.4 -36.43 2.5 -36.33 ;
        RECT 2.4 -37.96 2.5 -37.86 ;
        RECT 2.4 -38.315 2.5 -38.215 ;
        RECT 2.4 -39.305 2.5 -39.205 ;
        RECT 2.4 -39.66 2.5 -39.56 ;
        RECT 2.4 -41.19 2.5 -41.09 ;
        RECT 2.4 -41.545 2.5 -41.445 ;
        RECT 2.4 -42.535 2.5 -42.435 ;
        RECT 2.4 -42.89 2.5 -42.79 ;
        RECT 2.4 -44.42 2.5 -44.32 ;
        RECT 2.4 -44.775 2.5 -44.675 ;
        RECT 2.4 -45.765 2.5 -45.665 ;
        RECT 2.4 -46.12 2.5 -46.02 ;
        RECT 2.4 -47.65 2.5 -47.55 ;
        RECT 2.4 -48.005 2.5 -47.905 ;
        RECT 2.4 -48.995 2.5 -48.895 ;
        RECT 2.4 -49.35 2.5 -49.25 ;
        RECT 3.6 9.75 3.7 9.85 ;
        RECT 3.6 9.52 3.7 9.62 ;
        RECT 3.6 9.29 3.7 9.39 ;
        RECT 3.6 9.06 3.7 9.16 ;
        RECT 3.6 8.83 3.7 8.93 ;
        RECT 3.6 8.6 3.7 8.7 ;
        RECT 3.6 8.37 3.7 8.47 ;
        RECT 3.6 8.14 3.7 8.24 ;
        RECT 3.6 7.91 3.7 8.01 ;
        RECT 3.6 7.68 3.7 7.78 ;
        RECT 3.6 7.45 3.7 7.55 ;
        RECT 3.6 7.22 3.7 7.32 ;
        RECT 3.6 0.8 3.7 0.9 ;
        RECT 3.6 0.445 3.7 0.545 ;
        RECT 3.6 -0.545 3.7 -0.445 ;
        RECT 3.6 -0.9 3.7 -0.8 ;
        RECT 3.6 -2.43 3.7 -2.33 ;
        RECT 3.6 -2.785 3.7 -2.685 ;
        RECT 3.6 -3.775 3.7 -3.675 ;
        RECT 3.6 -4.13 3.7 -4.03 ;
        RECT 3.6 -5.66 3.7 -5.56 ;
        RECT 3.6 -6.015 3.7 -5.915 ;
        RECT 3.6 -7.005 3.7 -6.905 ;
        RECT 3.6 -7.36 3.7 -7.26 ;
        RECT 3.6 -8.89 3.7 -8.79 ;
        RECT 3.6 -9.245 3.7 -9.145 ;
        RECT 3.6 -10.235 3.7 -10.135 ;
        RECT 3.6 -10.59 3.7 -10.49 ;
        RECT 3.6 -12.12 3.7 -12.02 ;
        RECT 3.6 -12.475 3.7 -12.375 ;
        RECT 3.6 -13.465 3.7 -13.365 ;
        RECT 3.6 -13.82 3.7 -13.72 ;
        RECT 3.6 -15.35 3.7 -15.25 ;
        RECT 3.6 -15.705 3.7 -15.605 ;
        RECT 3.6 -16.695 3.7 -16.595 ;
        RECT 3.6 -17.05 3.7 -16.95 ;
        RECT 3.6 -18.58 3.7 -18.48 ;
        RECT 3.6 -18.935 3.7 -18.835 ;
        RECT 3.6 -19.925 3.7 -19.825 ;
        RECT 3.6 -20.28 3.7 -20.18 ;
        RECT 3.6 -21.81 3.7 -21.71 ;
        RECT 3.6 -22.165 3.7 -22.065 ;
        RECT 3.6 -23.155 3.7 -23.055 ;
        RECT 3.6 -23.51 3.7 -23.41 ;
        RECT 3.6 -25.04 3.7 -24.94 ;
        RECT 3.6 -25.395 3.7 -25.295 ;
        RECT 3.6 -26.385 3.7 -26.285 ;
        RECT 3.6 -26.74 3.7 -26.64 ;
        RECT 3.6 -28.27 3.7 -28.17 ;
        RECT 3.6 -28.625 3.7 -28.525 ;
        RECT 3.6 -29.615 3.7 -29.515 ;
        RECT 3.6 -29.97 3.7 -29.87 ;
        RECT 3.6 -31.5 3.7 -31.4 ;
        RECT 3.6 -31.855 3.7 -31.755 ;
        RECT 3.6 -32.845 3.7 -32.745 ;
        RECT 3.6 -33.2 3.7 -33.1 ;
        RECT 3.6 -34.73 3.7 -34.63 ;
        RECT 3.6 -35.085 3.7 -34.985 ;
        RECT 3.6 -36.075 3.7 -35.975 ;
        RECT 3.6 -36.43 3.7 -36.33 ;
        RECT 3.6 -37.96 3.7 -37.86 ;
        RECT 3.6 -38.315 3.7 -38.215 ;
        RECT 3.6 -39.305 3.7 -39.205 ;
        RECT 3.6 -39.66 3.7 -39.56 ;
        RECT 3.6 -41.19 3.7 -41.09 ;
        RECT 3.6 -41.545 3.7 -41.445 ;
        RECT 3.6 -42.535 3.7 -42.435 ;
        RECT 3.6 -42.89 3.7 -42.79 ;
        RECT 3.6 -44.42 3.7 -44.32 ;
        RECT 3.6 -44.775 3.7 -44.675 ;
        RECT 3.6 -45.765 3.7 -45.665 ;
        RECT 3.6 -46.12 3.7 -46.02 ;
        RECT 3.6 -47.65 3.7 -47.55 ;
        RECT 3.6 -48.005 3.7 -47.905 ;
        RECT 3.6 -48.995 3.7 -48.895 ;
        RECT 3.6 -49.35 3.7 -49.25 ;
        RECT 4.8 9.75 4.9 9.85 ;
        RECT 4.8 9.52 4.9 9.62 ;
        RECT 4.8 9.29 4.9 9.39 ;
        RECT 4.8 9.06 4.9 9.16 ;
        RECT 4.8 8.83 4.9 8.93 ;
        RECT 4.8 8.6 4.9 8.7 ;
        RECT 4.8 8.37 4.9 8.47 ;
        RECT 4.8 8.14 4.9 8.24 ;
        RECT 4.8 7.91 4.9 8.01 ;
        RECT 4.8 7.68 4.9 7.78 ;
        RECT 4.8 7.45 4.9 7.55 ;
        RECT 4.8 7.22 4.9 7.32 ;
        RECT 4.8 0.8 4.9 0.9 ;
        RECT 4.8 0.445 4.9 0.545 ;
        RECT 4.8 -0.545 4.9 -0.445 ;
        RECT 4.8 -0.9 4.9 -0.8 ;
        RECT 4.8 -2.43 4.9 -2.33 ;
        RECT 4.8 -2.785 4.9 -2.685 ;
        RECT 4.8 -3.775 4.9 -3.675 ;
        RECT 4.8 -4.13 4.9 -4.03 ;
        RECT 4.8 -5.66 4.9 -5.56 ;
        RECT 4.8 -6.015 4.9 -5.915 ;
        RECT 4.8 -7.005 4.9 -6.905 ;
        RECT 4.8 -7.36 4.9 -7.26 ;
        RECT 4.8 -8.89 4.9 -8.79 ;
        RECT 4.8 -9.245 4.9 -9.145 ;
        RECT 4.8 -10.235 4.9 -10.135 ;
        RECT 4.8 -10.59 4.9 -10.49 ;
        RECT 4.8 -12.12 4.9 -12.02 ;
        RECT 4.8 -12.475 4.9 -12.375 ;
        RECT 4.8 -13.465 4.9 -13.365 ;
        RECT 4.8 -13.82 4.9 -13.72 ;
        RECT 4.8 -15.35 4.9 -15.25 ;
        RECT 4.8 -15.705 4.9 -15.605 ;
        RECT 4.8 -16.695 4.9 -16.595 ;
        RECT 4.8 -17.05 4.9 -16.95 ;
        RECT 4.8 -18.58 4.9 -18.48 ;
        RECT 4.8 -18.935 4.9 -18.835 ;
        RECT 4.8 -19.925 4.9 -19.825 ;
        RECT 4.8 -20.28 4.9 -20.18 ;
        RECT 4.8 -21.81 4.9 -21.71 ;
        RECT 4.8 -22.165 4.9 -22.065 ;
        RECT 4.8 -23.155 4.9 -23.055 ;
        RECT 4.8 -23.51 4.9 -23.41 ;
        RECT 4.8 -25.04 4.9 -24.94 ;
        RECT 4.8 -25.395 4.9 -25.295 ;
        RECT 4.8 -26.385 4.9 -26.285 ;
        RECT 4.8 -26.74 4.9 -26.64 ;
        RECT 4.8 -28.27 4.9 -28.17 ;
        RECT 4.8 -28.625 4.9 -28.525 ;
        RECT 4.8 -29.615 4.9 -29.515 ;
        RECT 4.8 -29.97 4.9 -29.87 ;
        RECT 4.8 -31.5 4.9 -31.4 ;
        RECT 4.8 -31.855 4.9 -31.755 ;
        RECT 4.8 -32.845 4.9 -32.745 ;
        RECT 4.8 -33.2 4.9 -33.1 ;
        RECT 4.8 -34.73 4.9 -34.63 ;
        RECT 4.8 -35.085 4.9 -34.985 ;
        RECT 4.8 -36.075 4.9 -35.975 ;
        RECT 4.8 -36.43 4.9 -36.33 ;
        RECT 4.8 -37.96 4.9 -37.86 ;
        RECT 4.8 -38.315 4.9 -38.215 ;
        RECT 4.8 -39.305 4.9 -39.205 ;
        RECT 4.8 -39.66 4.9 -39.56 ;
        RECT 4.8 -41.19 4.9 -41.09 ;
        RECT 4.8 -41.545 4.9 -41.445 ;
        RECT 4.8 -42.535 4.9 -42.435 ;
        RECT 4.8 -42.89 4.9 -42.79 ;
        RECT 4.8 -44.42 4.9 -44.32 ;
        RECT 4.8 -44.775 4.9 -44.675 ;
        RECT 4.8 -45.765 4.9 -45.665 ;
        RECT 4.8 -46.12 4.9 -46.02 ;
        RECT 4.8 -47.65 4.9 -47.55 ;
        RECT 4.8 -48.005 4.9 -47.905 ;
        RECT 4.8 -48.995 4.9 -48.895 ;
        RECT 4.8 -49.35 4.9 -49.25 ;
        RECT 6 9.75 6.1 9.85 ;
        RECT 6 9.52 6.1 9.62 ;
        RECT 6 9.29 6.1 9.39 ;
        RECT 6 9.06 6.1 9.16 ;
        RECT 6 8.83 6.1 8.93 ;
        RECT 6 8.6 6.1 8.7 ;
        RECT 6 8.37 6.1 8.47 ;
        RECT 6 8.14 6.1 8.24 ;
        RECT 6 7.91 6.1 8.01 ;
        RECT 6 7.68 6.1 7.78 ;
        RECT 6 7.45 6.1 7.55 ;
        RECT 6 7.22 6.1 7.32 ;
        RECT 6 0.8 6.1 0.9 ;
        RECT 6 0.445 6.1 0.545 ;
        RECT 6 -0.545 6.1 -0.445 ;
        RECT 6 -0.9 6.1 -0.8 ;
        RECT 6 -2.43 6.1 -2.33 ;
        RECT 6 -2.785 6.1 -2.685 ;
        RECT 6 -3.775 6.1 -3.675 ;
        RECT 6 -4.13 6.1 -4.03 ;
        RECT 6 -5.66 6.1 -5.56 ;
        RECT 6 -6.015 6.1 -5.915 ;
        RECT 6 -7.005 6.1 -6.905 ;
        RECT 6 -7.36 6.1 -7.26 ;
        RECT 6 -8.89 6.1 -8.79 ;
        RECT 6 -9.245 6.1 -9.145 ;
        RECT 6 -10.235 6.1 -10.135 ;
        RECT 6 -10.59 6.1 -10.49 ;
        RECT 6 -12.12 6.1 -12.02 ;
        RECT 6 -12.475 6.1 -12.375 ;
        RECT 6 -13.465 6.1 -13.365 ;
        RECT 6 -13.82 6.1 -13.72 ;
        RECT 6 -15.35 6.1 -15.25 ;
        RECT 6 -15.705 6.1 -15.605 ;
        RECT 6 -16.695 6.1 -16.595 ;
        RECT 6 -17.05 6.1 -16.95 ;
        RECT 6 -18.58 6.1 -18.48 ;
        RECT 6 -18.935 6.1 -18.835 ;
        RECT 6 -19.925 6.1 -19.825 ;
        RECT 6 -20.28 6.1 -20.18 ;
        RECT 6 -21.81 6.1 -21.71 ;
        RECT 6 -22.165 6.1 -22.065 ;
        RECT 6 -23.155 6.1 -23.055 ;
        RECT 6 -23.51 6.1 -23.41 ;
        RECT 6 -25.04 6.1 -24.94 ;
        RECT 6 -25.395 6.1 -25.295 ;
        RECT 6 -26.385 6.1 -26.285 ;
        RECT 6 -26.74 6.1 -26.64 ;
        RECT 6 -28.27 6.1 -28.17 ;
        RECT 6 -28.625 6.1 -28.525 ;
        RECT 6 -29.615 6.1 -29.515 ;
        RECT 6 -29.97 6.1 -29.87 ;
        RECT 6 -31.5 6.1 -31.4 ;
        RECT 6 -31.855 6.1 -31.755 ;
        RECT 6 -32.845 6.1 -32.745 ;
        RECT 6 -33.2 6.1 -33.1 ;
        RECT 6 -34.73 6.1 -34.63 ;
        RECT 6 -35.085 6.1 -34.985 ;
        RECT 6 -36.075 6.1 -35.975 ;
        RECT 6 -36.43 6.1 -36.33 ;
        RECT 6 -37.96 6.1 -37.86 ;
        RECT 6 -38.315 6.1 -38.215 ;
        RECT 6 -39.305 6.1 -39.205 ;
        RECT 6 -39.66 6.1 -39.56 ;
        RECT 6 -41.19 6.1 -41.09 ;
        RECT 6 -41.545 6.1 -41.445 ;
        RECT 6 -42.535 6.1 -42.435 ;
        RECT 6 -42.89 6.1 -42.79 ;
        RECT 6 -44.42 6.1 -44.32 ;
        RECT 6 -44.775 6.1 -44.675 ;
        RECT 6 -45.765 6.1 -45.665 ;
        RECT 6 -46.12 6.1 -46.02 ;
        RECT 6 -47.65 6.1 -47.55 ;
        RECT 6 -48.005 6.1 -47.905 ;
        RECT 6 -48.995 6.1 -48.895 ;
        RECT 6 -49.35 6.1 -49.25 ;
        RECT 7.2 9.75 7.3 9.85 ;
        RECT 7.2 9.52 7.3 9.62 ;
        RECT 7.2 9.29 7.3 9.39 ;
        RECT 7.2 9.06 7.3 9.16 ;
        RECT 7.2 8.83 7.3 8.93 ;
        RECT 7.2 8.6 7.3 8.7 ;
        RECT 7.2 8.37 7.3 8.47 ;
        RECT 7.2 8.14 7.3 8.24 ;
        RECT 7.2 7.91 7.3 8.01 ;
        RECT 7.2 7.68 7.3 7.78 ;
        RECT 7.2 7.45 7.3 7.55 ;
        RECT 7.2 7.22 7.3 7.32 ;
        RECT 7.2 0.8 7.3 0.9 ;
        RECT 7.2 0.445 7.3 0.545 ;
        RECT 7.2 -0.545 7.3 -0.445 ;
        RECT 7.2 -0.9 7.3 -0.8 ;
        RECT 7.2 -2.43 7.3 -2.33 ;
        RECT 7.2 -2.785 7.3 -2.685 ;
        RECT 7.2 -3.775 7.3 -3.675 ;
        RECT 7.2 -4.13 7.3 -4.03 ;
        RECT 7.2 -5.66 7.3 -5.56 ;
        RECT 7.2 -6.015 7.3 -5.915 ;
        RECT 7.2 -7.005 7.3 -6.905 ;
        RECT 7.2 -7.36 7.3 -7.26 ;
        RECT 7.2 -8.89 7.3 -8.79 ;
        RECT 7.2 -9.245 7.3 -9.145 ;
        RECT 7.2 -10.235 7.3 -10.135 ;
        RECT 7.2 -10.59 7.3 -10.49 ;
        RECT 7.2 -12.12 7.3 -12.02 ;
        RECT 7.2 -12.475 7.3 -12.375 ;
        RECT 7.2 -13.465 7.3 -13.365 ;
        RECT 7.2 -13.82 7.3 -13.72 ;
        RECT 7.2 -15.35 7.3 -15.25 ;
        RECT 7.2 -15.705 7.3 -15.605 ;
        RECT 7.2 -16.695 7.3 -16.595 ;
        RECT 7.2 -17.05 7.3 -16.95 ;
        RECT 7.2 -18.58 7.3 -18.48 ;
        RECT 7.2 -18.935 7.3 -18.835 ;
        RECT 7.2 -19.925 7.3 -19.825 ;
        RECT 7.2 -20.28 7.3 -20.18 ;
        RECT 7.2 -21.81 7.3 -21.71 ;
        RECT 7.2 -22.165 7.3 -22.065 ;
        RECT 7.2 -23.155 7.3 -23.055 ;
        RECT 7.2 -23.51 7.3 -23.41 ;
        RECT 7.2 -25.04 7.3 -24.94 ;
        RECT 7.2 -25.395 7.3 -25.295 ;
        RECT 7.2 -26.385 7.3 -26.285 ;
        RECT 7.2 -26.74 7.3 -26.64 ;
        RECT 7.2 -28.27 7.3 -28.17 ;
        RECT 7.2 -28.625 7.3 -28.525 ;
        RECT 7.2 -29.615 7.3 -29.515 ;
        RECT 7.2 -29.97 7.3 -29.87 ;
        RECT 7.2 -31.5 7.3 -31.4 ;
        RECT 7.2 -31.855 7.3 -31.755 ;
        RECT 7.2 -32.845 7.3 -32.745 ;
        RECT 7.2 -33.2 7.3 -33.1 ;
        RECT 7.2 -34.73 7.3 -34.63 ;
        RECT 7.2 -35.085 7.3 -34.985 ;
        RECT 7.2 -36.075 7.3 -35.975 ;
        RECT 7.2 -36.43 7.3 -36.33 ;
        RECT 7.2 -37.96 7.3 -37.86 ;
        RECT 7.2 -38.315 7.3 -38.215 ;
        RECT 7.2 -39.305 7.3 -39.205 ;
        RECT 7.2 -39.66 7.3 -39.56 ;
        RECT 7.2 -41.19 7.3 -41.09 ;
        RECT 7.2 -41.545 7.3 -41.445 ;
        RECT 7.2 -42.535 7.3 -42.435 ;
        RECT 7.2 -42.89 7.3 -42.79 ;
        RECT 7.2 -44.42 7.3 -44.32 ;
        RECT 7.2 -44.775 7.3 -44.675 ;
        RECT 7.2 -45.765 7.3 -45.665 ;
        RECT 7.2 -46.12 7.3 -46.02 ;
        RECT 7.2 -47.65 7.3 -47.55 ;
        RECT 7.2 -48.005 7.3 -47.905 ;
        RECT 7.2 -48.995 7.3 -48.895 ;
        RECT 7.2 -49.35 7.3 -49.25 ;
        RECT 8.4 9.75 8.5 9.85 ;
        RECT 8.4 9.52 8.5 9.62 ;
        RECT 8.4 9.29 8.5 9.39 ;
        RECT 8.4 9.06 8.5 9.16 ;
        RECT 8.4 8.83 8.5 8.93 ;
        RECT 8.4 8.6 8.5 8.7 ;
        RECT 8.4 8.37 8.5 8.47 ;
        RECT 8.4 8.14 8.5 8.24 ;
        RECT 8.4 7.91 8.5 8.01 ;
        RECT 8.4 7.68 8.5 7.78 ;
        RECT 8.4 7.45 8.5 7.55 ;
        RECT 8.4 7.22 8.5 7.32 ;
        RECT 8.4 0.8 8.5 0.9 ;
        RECT 8.4 0.445 8.5 0.545 ;
        RECT 8.4 -0.545 8.5 -0.445 ;
        RECT 8.4 -0.9 8.5 -0.8 ;
        RECT 8.4 -2.43 8.5 -2.33 ;
        RECT 8.4 -2.785 8.5 -2.685 ;
        RECT 8.4 -3.775 8.5 -3.675 ;
        RECT 8.4 -4.13 8.5 -4.03 ;
        RECT 8.4 -5.66 8.5 -5.56 ;
        RECT 8.4 -6.015 8.5 -5.915 ;
        RECT 8.4 -7.005 8.5 -6.905 ;
        RECT 8.4 -7.36 8.5 -7.26 ;
        RECT 8.4 -8.89 8.5 -8.79 ;
        RECT 8.4 -9.245 8.5 -9.145 ;
        RECT 8.4 -10.235 8.5 -10.135 ;
        RECT 8.4 -10.59 8.5 -10.49 ;
        RECT 8.4 -12.12 8.5 -12.02 ;
        RECT 8.4 -12.475 8.5 -12.375 ;
        RECT 8.4 -13.465 8.5 -13.365 ;
        RECT 8.4 -13.82 8.5 -13.72 ;
        RECT 8.4 -15.35 8.5 -15.25 ;
        RECT 8.4 -15.705 8.5 -15.605 ;
        RECT 8.4 -16.695 8.5 -16.595 ;
        RECT 8.4 -17.05 8.5 -16.95 ;
        RECT 8.4 -18.58 8.5 -18.48 ;
        RECT 8.4 -18.935 8.5 -18.835 ;
        RECT 8.4 -19.925 8.5 -19.825 ;
        RECT 8.4 -20.28 8.5 -20.18 ;
        RECT 8.4 -21.81 8.5 -21.71 ;
        RECT 8.4 -22.165 8.5 -22.065 ;
        RECT 8.4 -23.155 8.5 -23.055 ;
        RECT 8.4 -23.51 8.5 -23.41 ;
        RECT 8.4 -25.04 8.5 -24.94 ;
        RECT 8.4 -25.395 8.5 -25.295 ;
        RECT 8.4 -26.385 8.5 -26.285 ;
        RECT 8.4 -26.74 8.5 -26.64 ;
        RECT 8.4 -28.27 8.5 -28.17 ;
        RECT 8.4 -28.625 8.5 -28.525 ;
        RECT 8.4 -29.615 8.5 -29.515 ;
        RECT 8.4 -29.97 8.5 -29.87 ;
        RECT 8.4 -31.5 8.5 -31.4 ;
        RECT 8.4 -31.855 8.5 -31.755 ;
        RECT 8.4 -32.845 8.5 -32.745 ;
        RECT 8.4 -33.2 8.5 -33.1 ;
        RECT 8.4 -34.73 8.5 -34.63 ;
        RECT 8.4 -35.085 8.5 -34.985 ;
        RECT 8.4 -36.075 8.5 -35.975 ;
        RECT 8.4 -36.43 8.5 -36.33 ;
        RECT 8.4 -37.96 8.5 -37.86 ;
        RECT 8.4 -38.315 8.5 -38.215 ;
        RECT 8.4 -39.305 8.5 -39.205 ;
        RECT 8.4 -39.66 8.5 -39.56 ;
        RECT 8.4 -41.19 8.5 -41.09 ;
        RECT 8.4 -41.545 8.5 -41.445 ;
        RECT 8.4 -42.535 8.5 -42.435 ;
        RECT 8.4 -42.89 8.5 -42.79 ;
        RECT 8.4 -44.42 8.5 -44.32 ;
        RECT 8.4 -44.775 8.5 -44.675 ;
        RECT 8.4 -45.765 8.5 -45.665 ;
        RECT 8.4 -46.12 8.5 -46.02 ;
        RECT 8.4 -47.65 8.5 -47.55 ;
        RECT 8.4 -48.005 8.5 -47.905 ;
        RECT 8.4 -48.995 8.5 -48.895 ;
        RECT 8.4 -49.35 8.5 -49.25 ;
        RECT 9.6 9.75 9.7 9.85 ;
        RECT 9.6 9.52 9.7 9.62 ;
        RECT 9.6 9.29 9.7 9.39 ;
        RECT 9.6 9.06 9.7 9.16 ;
        RECT 9.6 8.83 9.7 8.93 ;
        RECT 9.6 8.6 9.7 8.7 ;
        RECT 9.6 8.37 9.7 8.47 ;
        RECT 9.6 8.14 9.7 8.24 ;
        RECT 9.6 7.91 9.7 8.01 ;
        RECT 9.6 7.68 9.7 7.78 ;
        RECT 9.6 7.45 9.7 7.55 ;
        RECT 9.6 7.22 9.7 7.32 ;
        RECT 9.6 0.8 9.7 0.9 ;
        RECT 9.6 0.445 9.7 0.545 ;
        RECT 9.6 -0.545 9.7 -0.445 ;
        RECT 9.6 -0.9 9.7 -0.8 ;
        RECT 9.6 -2.43 9.7 -2.33 ;
        RECT 9.6 -2.785 9.7 -2.685 ;
        RECT 9.6 -3.775 9.7 -3.675 ;
        RECT 9.6 -4.13 9.7 -4.03 ;
        RECT 9.6 -5.66 9.7 -5.56 ;
        RECT 9.6 -6.015 9.7 -5.915 ;
        RECT 9.6 -7.005 9.7 -6.905 ;
        RECT 9.6 -7.36 9.7 -7.26 ;
        RECT 9.6 -8.89 9.7 -8.79 ;
        RECT 9.6 -9.245 9.7 -9.145 ;
        RECT 9.6 -10.235 9.7 -10.135 ;
        RECT 9.6 -10.59 9.7 -10.49 ;
        RECT 9.6 -12.12 9.7 -12.02 ;
        RECT 9.6 -12.475 9.7 -12.375 ;
        RECT 9.6 -13.465 9.7 -13.365 ;
        RECT 9.6 -13.82 9.7 -13.72 ;
        RECT 9.6 -15.35 9.7 -15.25 ;
        RECT 9.6 -15.705 9.7 -15.605 ;
        RECT 9.6 -16.695 9.7 -16.595 ;
        RECT 9.6 -17.05 9.7 -16.95 ;
        RECT 9.6 -18.58 9.7 -18.48 ;
        RECT 9.6 -18.935 9.7 -18.835 ;
        RECT 9.6 -19.925 9.7 -19.825 ;
        RECT 9.6 -20.28 9.7 -20.18 ;
        RECT 9.6 -21.81 9.7 -21.71 ;
        RECT 9.6 -22.165 9.7 -22.065 ;
        RECT 9.6 -23.155 9.7 -23.055 ;
        RECT 9.6 -23.51 9.7 -23.41 ;
        RECT 9.6 -25.04 9.7 -24.94 ;
        RECT 9.6 -25.395 9.7 -25.295 ;
        RECT 9.6 -26.385 9.7 -26.285 ;
        RECT 9.6 -26.74 9.7 -26.64 ;
        RECT 9.6 -28.27 9.7 -28.17 ;
        RECT 9.6 -28.625 9.7 -28.525 ;
        RECT 9.6 -29.615 9.7 -29.515 ;
        RECT 9.6 -29.97 9.7 -29.87 ;
        RECT 9.6 -31.5 9.7 -31.4 ;
        RECT 9.6 -31.855 9.7 -31.755 ;
        RECT 9.6 -32.845 9.7 -32.745 ;
        RECT 9.6 -33.2 9.7 -33.1 ;
        RECT 9.6 -34.73 9.7 -34.63 ;
        RECT 9.6 -35.085 9.7 -34.985 ;
        RECT 9.6 -36.075 9.7 -35.975 ;
        RECT 9.6 -36.43 9.7 -36.33 ;
        RECT 9.6 -37.96 9.7 -37.86 ;
        RECT 9.6 -38.315 9.7 -38.215 ;
        RECT 9.6 -39.305 9.7 -39.205 ;
        RECT 9.6 -39.66 9.7 -39.56 ;
        RECT 9.6 -41.19 9.7 -41.09 ;
        RECT 9.6 -41.545 9.7 -41.445 ;
        RECT 9.6 -42.535 9.7 -42.435 ;
        RECT 9.6 -42.89 9.7 -42.79 ;
        RECT 9.6 -44.42 9.7 -44.32 ;
        RECT 9.6 -44.775 9.7 -44.675 ;
        RECT 9.6 -45.765 9.7 -45.665 ;
        RECT 9.6 -46.12 9.7 -46.02 ;
        RECT 9.6 -47.65 9.7 -47.55 ;
        RECT 9.6 -48.005 9.7 -47.905 ;
        RECT 9.6 -48.995 9.7 -48.895 ;
        RECT 9.6 -49.35 9.7 -49.25 ;
        RECT 10.8 9.75 10.9 9.85 ;
        RECT 10.8 9.52 10.9 9.62 ;
        RECT 10.8 9.29 10.9 9.39 ;
        RECT 10.8 9.06 10.9 9.16 ;
        RECT 10.8 8.83 10.9 8.93 ;
        RECT 10.8 8.6 10.9 8.7 ;
        RECT 10.8 8.37 10.9 8.47 ;
        RECT 10.8 8.14 10.9 8.24 ;
        RECT 10.8 7.91 10.9 8.01 ;
        RECT 10.8 7.68 10.9 7.78 ;
        RECT 10.8 7.45 10.9 7.55 ;
        RECT 10.8 7.22 10.9 7.32 ;
        RECT 10.8 0.8 10.9 0.9 ;
        RECT 10.8 0.445 10.9 0.545 ;
        RECT 10.8 -0.545 10.9 -0.445 ;
        RECT 10.8 -0.9 10.9 -0.8 ;
        RECT 10.8 -2.43 10.9 -2.33 ;
        RECT 10.8 -2.785 10.9 -2.685 ;
        RECT 10.8 -3.775 10.9 -3.675 ;
        RECT 10.8 -4.13 10.9 -4.03 ;
        RECT 10.8 -5.66 10.9 -5.56 ;
        RECT 10.8 -6.015 10.9 -5.915 ;
        RECT 10.8 -7.005 10.9 -6.905 ;
        RECT 10.8 -7.36 10.9 -7.26 ;
        RECT 10.8 -8.89 10.9 -8.79 ;
        RECT 10.8 -9.245 10.9 -9.145 ;
        RECT 10.8 -10.235 10.9 -10.135 ;
        RECT 10.8 -10.59 10.9 -10.49 ;
        RECT 10.8 -12.12 10.9 -12.02 ;
        RECT 10.8 -12.475 10.9 -12.375 ;
        RECT 10.8 -13.465 10.9 -13.365 ;
        RECT 10.8 -13.82 10.9 -13.72 ;
        RECT 10.8 -15.35 10.9 -15.25 ;
        RECT 10.8 -15.705 10.9 -15.605 ;
        RECT 10.8 -16.695 10.9 -16.595 ;
        RECT 10.8 -17.05 10.9 -16.95 ;
        RECT 10.8 -18.58 10.9 -18.48 ;
        RECT 10.8 -18.935 10.9 -18.835 ;
        RECT 10.8 -19.925 10.9 -19.825 ;
        RECT 10.8 -20.28 10.9 -20.18 ;
        RECT 10.8 -21.81 10.9 -21.71 ;
        RECT 10.8 -22.165 10.9 -22.065 ;
        RECT 10.8 -23.155 10.9 -23.055 ;
        RECT 10.8 -23.51 10.9 -23.41 ;
        RECT 10.8 -25.04 10.9 -24.94 ;
        RECT 10.8 -25.395 10.9 -25.295 ;
        RECT 10.8 -26.385 10.9 -26.285 ;
        RECT 10.8 -26.74 10.9 -26.64 ;
        RECT 10.8 -28.27 10.9 -28.17 ;
        RECT 10.8 -28.625 10.9 -28.525 ;
        RECT 10.8 -29.615 10.9 -29.515 ;
        RECT 10.8 -29.97 10.9 -29.87 ;
        RECT 10.8 -31.5 10.9 -31.4 ;
        RECT 10.8 -31.855 10.9 -31.755 ;
        RECT 10.8 -32.845 10.9 -32.745 ;
        RECT 10.8 -33.2 10.9 -33.1 ;
        RECT 10.8 -34.73 10.9 -34.63 ;
        RECT 10.8 -35.085 10.9 -34.985 ;
        RECT 10.8 -36.075 10.9 -35.975 ;
        RECT 10.8 -36.43 10.9 -36.33 ;
        RECT 10.8 -37.96 10.9 -37.86 ;
        RECT 10.8 -38.315 10.9 -38.215 ;
        RECT 10.8 -39.305 10.9 -39.205 ;
        RECT 10.8 -39.66 10.9 -39.56 ;
        RECT 10.8 -41.19 10.9 -41.09 ;
        RECT 10.8 -41.545 10.9 -41.445 ;
        RECT 10.8 -42.535 10.9 -42.435 ;
        RECT 10.8 -42.89 10.9 -42.79 ;
        RECT 10.8 -44.42 10.9 -44.32 ;
        RECT 10.8 -44.775 10.9 -44.675 ;
        RECT 10.8 -45.765 10.9 -45.665 ;
        RECT 10.8 -46.12 10.9 -46.02 ;
        RECT 10.8 -47.65 10.9 -47.55 ;
        RECT 10.8 -48.005 10.9 -47.905 ;
        RECT 10.8 -48.995 10.9 -48.895 ;
        RECT 10.8 -49.35 10.9 -49.25 ;
        RECT 12 9.75 12.1 9.85 ;
        RECT 12 9.52 12.1 9.62 ;
        RECT 12 9.29 12.1 9.39 ;
        RECT 12 9.06 12.1 9.16 ;
        RECT 12 8.83 12.1 8.93 ;
        RECT 12 8.6 12.1 8.7 ;
        RECT 12 8.37 12.1 8.47 ;
        RECT 12 8.14 12.1 8.24 ;
        RECT 12 7.91 12.1 8.01 ;
        RECT 12 7.68 12.1 7.78 ;
        RECT 12 7.45 12.1 7.55 ;
        RECT 12 7.22 12.1 7.32 ;
        RECT 12 0.8 12.1 0.9 ;
        RECT 12 0.445 12.1 0.545 ;
        RECT 12 -0.545 12.1 -0.445 ;
        RECT 12 -0.9 12.1 -0.8 ;
        RECT 12 -2.43 12.1 -2.33 ;
        RECT 12 -2.785 12.1 -2.685 ;
        RECT 12 -3.775 12.1 -3.675 ;
        RECT 12 -4.13 12.1 -4.03 ;
        RECT 12 -5.66 12.1 -5.56 ;
        RECT 12 -6.015 12.1 -5.915 ;
        RECT 12 -7.005 12.1 -6.905 ;
        RECT 12 -7.36 12.1 -7.26 ;
        RECT 12 -8.89 12.1 -8.79 ;
        RECT 12 -9.245 12.1 -9.145 ;
        RECT 12 -10.235 12.1 -10.135 ;
        RECT 12 -10.59 12.1 -10.49 ;
        RECT 12 -12.12 12.1 -12.02 ;
        RECT 12 -12.475 12.1 -12.375 ;
        RECT 12 -13.465 12.1 -13.365 ;
        RECT 12 -13.82 12.1 -13.72 ;
        RECT 12 -15.35 12.1 -15.25 ;
        RECT 12 -15.705 12.1 -15.605 ;
        RECT 12 -16.695 12.1 -16.595 ;
        RECT 12 -17.05 12.1 -16.95 ;
        RECT 12 -18.58 12.1 -18.48 ;
        RECT 12 -18.935 12.1 -18.835 ;
        RECT 12 -19.925 12.1 -19.825 ;
        RECT 12 -20.28 12.1 -20.18 ;
        RECT 12 -21.81 12.1 -21.71 ;
        RECT 12 -22.165 12.1 -22.065 ;
        RECT 12 -23.155 12.1 -23.055 ;
        RECT 12 -23.51 12.1 -23.41 ;
        RECT 12 -25.04 12.1 -24.94 ;
        RECT 12 -25.395 12.1 -25.295 ;
        RECT 12 -26.385 12.1 -26.285 ;
        RECT 12 -26.74 12.1 -26.64 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INPUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER M2 ;
        RECT 40.265 -68.685 41.265 5.175 ;
        RECT -31.525 -68.925 -30.525 5.645 ;
      LAYER M1 ;
        RECT -33.525 -68.685 43.265 -65.965 ;
        RECT 0.01 -61.145 41.265 -60.785 ;
        RECT 38.005 -61.145 38.105 -60.095 ;
        RECT 37.445 -61.145 37.545 -60.095 ;
        RECT 36.855 -61.145 36.955 -60.095 ;
        RECT 36.295 -61.145 36.395 -60.095 ;
        RECT 35.985 -61.145 36.085 -60.095 ;
        RECT 35.83 -61.595 35.93 -60.785 ;
        RECT 35.425 -61.145 35.525 -60.095 ;
        RECT 35.24 -61.595 35.34 -60.785 ;
        RECT 34.835 -61.145 34.935 -60.095 ;
        RECT 34.275 -61.145 34.375 -60.095 ;
        RECT 33.685 -61.145 33.785 -60.095 ;
        RECT 33.205 -61.145 33.305 -60.095 ;
        RECT 32.645 -61.145 32.745 -60.095 ;
        RECT 32.055 -61.145 32.155 -60.095 ;
        RECT 31.495 -61.145 31.595 -60.095 ;
        RECT 31.185 -61.145 31.285 -60.095 ;
        RECT 31.03 -61.595 31.13 -60.785 ;
        RECT 30.625 -61.145 30.725 -60.095 ;
        RECT 30.44 -61.595 30.54 -60.785 ;
        RECT 30.035 -61.145 30.135 -60.095 ;
        RECT 29.475 -61.145 29.575 -60.095 ;
        RECT 28.885 -61.145 28.985 -60.095 ;
        RECT 28.405 -61.145 28.505 -60.095 ;
        RECT 27.845 -61.145 27.945 -60.095 ;
        RECT 27.255 -61.145 27.355 -60.095 ;
        RECT 26.695 -61.145 26.795 -60.095 ;
        RECT 26.385 -61.145 26.485 -60.095 ;
        RECT 26.23 -61.595 26.33 -60.785 ;
        RECT 25.825 -61.145 25.925 -60.095 ;
        RECT 25.64 -61.595 25.74 -60.785 ;
        RECT 25.235 -61.145 25.335 -60.095 ;
        RECT 24.675 -61.145 24.775 -60.095 ;
        RECT 24.085 -61.145 24.185 -60.095 ;
        RECT 23.605 -61.145 23.705 -60.095 ;
        RECT 23.045 -61.145 23.145 -60.095 ;
        RECT 22.455 -61.145 22.555 -60.095 ;
        RECT 21.895 -61.145 21.995 -60.095 ;
        RECT 21.585 -61.145 21.685 -60.095 ;
        RECT 21.43 -61.595 21.53 -60.785 ;
        RECT 21.025 -61.145 21.125 -60.095 ;
        RECT 20.84 -61.595 20.94 -60.785 ;
        RECT 20.435 -61.145 20.535 -60.095 ;
        RECT 19.875 -61.145 19.975 -60.095 ;
        RECT 19.285 -61.145 19.385 -60.095 ;
        RECT 18.805 -61.145 18.905 -60.095 ;
        RECT 18.245 -61.145 18.345 -60.095 ;
        RECT 17.655 -61.145 17.755 -60.095 ;
        RECT 17.095 -61.145 17.195 -60.095 ;
        RECT 16.785 -61.145 16.885 -60.095 ;
        RECT 16.63 -61.595 16.73 -60.785 ;
        RECT 16.225 -61.145 16.325 -60.095 ;
        RECT 16.04 -61.595 16.14 -60.785 ;
        RECT 15.635 -61.145 15.735 -60.095 ;
        RECT 15.075 -61.145 15.175 -60.095 ;
        RECT 14.485 -61.145 14.585 -60.095 ;
        RECT 14.005 -61.145 14.105 -60.095 ;
        RECT 13.445 -61.145 13.545 -60.095 ;
        RECT 12.855 -61.145 12.955 -60.095 ;
        RECT 12.295 -61.145 12.395 -60.095 ;
        RECT 11.985 -61.145 12.085 -60.095 ;
        RECT 11.83 -61.595 11.93 -60.785 ;
        RECT 11.425 -61.145 11.525 -60.095 ;
        RECT 11.24 -61.595 11.34 -60.785 ;
        RECT 10.835 -61.145 10.935 -60.095 ;
        RECT 10.275 -61.145 10.375 -60.095 ;
        RECT 9.685 -61.145 9.785 -60.095 ;
        RECT 9.205 -61.145 9.305 -60.095 ;
        RECT 8.645 -61.145 8.745 -60.095 ;
        RECT 8.055 -61.145 8.155 -60.095 ;
        RECT 7.495 -61.145 7.595 -60.095 ;
        RECT 7.185 -61.145 7.285 -60.095 ;
        RECT 7.03 -61.595 7.13 -60.785 ;
        RECT 6.625 -61.145 6.725 -60.095 ;
        RECT 6.44 -61.595 6.54 -60.785 ;
        RECT 6.035 -61.145 6.135 -60.095 ;
        RECT 5.475 -61.145 5.575 -60.095 ;
        RECT 4.885 -61.145 4.985 -60.095 ;
        RECT 4.405 -61.145 4.505 -60.095 ;
        RECT 3.845 -61.145 3.945 -60.095 ;
        RECT 3.255 -61.145 3.355 -60.095 ;
        RECT 2.695 -61.145 2.795 -60.095 ;
        RECT 2.385 -61.145 2.485 -60.095 ;
        RECT 2.23 -61.595 2.33 -60.785 ;
        RECT 1.825 -61.145 1.925 -60.095 ;
        RECT 1.64 -61.595 1.74 -60.785 ;
        RECT 1.235 -61.145 1.335 -60.095 ;
        RECT 0.675 -61.145 0.775 -60.095 ;
        RECT 0.085 -61.145 0.185 -60.095 ;
        RECT -0.055 -50.125 41.265 -50.005 ;
        RECT 38.4 -50.125 38.5 -49.66 ;
        RECT 37.2 -50.125 37.3 -49.66 ;
        RECT 36 -50.125 36.1 -49.66 ;
        RECT 34.8 -50.125 34.9 -49.66 ;
        RECT 33.6 -50.125 33.7 -49.66 ;
        RECT 32.4 -50.125 32.5 -49.66 ;
        RECT 31.2 -50.125 31.3 -49.66 ;
        RECT 30 -50.125 30.1 -49.66 ;
        RECT 28.8 -50.125 28.9 -49.66 ;
        RECT 27.6 -50.125 27.7 -49.66 ;
        RECT 26.4 -50.125 26.5 -49.66 ;
        RECT 25.2 -50.125 25.3 -49.66 ;
        RECT 24 -50.125 24.1 -49.66 ;
        RECT 22.8 -50.125 22.9 -49.66 ;
        RECT 21.6 -50.125 21.7 -49.66 ;
        RECT 20.4 -50.125 20.5 -49.66 ;
        RECT 19.2 -50.125 19.3 -49.66 ;
        RECT 18 -50.125 18.1 -49.66 ;
        RECT 16.8 -50.125 16.9 -49.66 ;
        RECT 15.6 -50.125 15.7 -49.66 ;
        RECT 14.4 -50.125 14.5 -49.66 ;
        RECT 13.2 -50.125 13.3 -49.66 ;
        RECT 12 -50.125 12.1 -49.66 ;
        RECT 10.8 -50.125 10.9 -49.66 ;
        RECT 9.6 -50.125 9.7 -49.66 ;
        RECT 8.4 -50.125 8.5 -49.66 ;
        RECT 7.2 -50.125 7.3 -49.66 ;
        RECT 6 -50.125 6.1 -49.66 ;
        RECT 4.8 -50.125 4.9 -49.66 ;
        RECT 3.6 -50.125 3.7 -49.66 ;
        RECT 2.4 -50.125 2.5 -49.66 ;
        RECT 1.2 -50.125 1.3 -49.66 ;
        RECT 0 -50.125 0.1 -49.66 ;
        RECT -0.055 -46.895 41.265 -46.775 ;
        RECT 38.4 -47.24 38.5 -46.43 ;
        RECT 37.2 -47.24 37.3 -46.43 ;
        RECT 36 -47.24 36.1 -46.43 ;
        RECT 34.8 -47.24 34.9 -46.43 ;
        RECT 33.6 -47.24 33.7 -46.43 ;
        RECT 32.4 -47.24 32.5 -46.43 ;
        RECT 31.2 -47.24 31.3 -46.43 ;
        RECT 30 -47.24 30.1 -46.43 ;
        RECT 28.8 -47.24 28.9 -46.43 ;
        RECT 27.6 -47.24 27.7 -46.43 ;
        RECT 26.4 -47.24 26.5 -46.43 ;
        RECT 25.2 -47.24 25.3 -46.43 ;
        RECT 24 -47.24 24.1 -46.43 ;
        RECT 22.8 -47.24 22.9 -46.43 ;
        RECT 21.6 -47.24 21.7 -46.43 ;
        RECT 20.4 -47.24 20.5 -46.43 ;
        RECT 19.2 -47.24 19.3 -46.43 ;
        RECT 18 -47.24 18.1 -46.43 ;
        RECT 16.8 -47.24 16.9 -46.43 ;
        RECT 15.6 -47.24 15.7 -46.43 ;
        RECT 14.4 -47.24 14.5 -46.43 ;
        RECT 13.2 -47.24 13.3 -46.43 ;
        RECT 12 -47.24 12.1 -46.43 ;
        RECT 10.8 -47.24 10.9 -46.43 ;
        RECT 9.6 -47.24 9.7 -46.43 ;
        RECT 8.4 -47.24 8.5 -46.43 ;
        RECT 7.2 -47.24 7.3 -46.43 ;
        RECT 6 -47.24 6.1 -46.43 ;
        RECT 4.8 -47.24 4.9 -46.43 ;
        RECT 3.6 -47.24 3.7 -46.43 ;
        RECT 2.4 -47.24 2.5 -46.43 ;
        RECT 1.2 -47.24 1.3 -46.43 ;
        RECT 0 -47.24 0.1 -46.43 ;
        RECT -0.055 -43.665 41.265 -43.545 ;
        RECT 38.4 -44.01 38.5 -43.2 ;
        RECT 37.2 -44.01 37.3 -43.2 ;
        RECT 36 -44.01 36.1 -43.2 ;
        RECT 34.8 -44.01 34.9 -43.2 ;
        RECT 33.6 -44.01 33.7 -43.2 ;
        RECT 32.4 -44.01 32.5 -43.2 ;
        RECT 31.2 -44.01 31.3 -43.2 ;
        RECT 30 -44.01 30.1 -43.2 ;
        RECT 28.8 -44.01 28.9 -43.2 ;
        RECT 27.6 -44.01 27.7 -43.2 ;
        RECT 26.4 -44.01 26.5 -43.2 ;
        RECT 25.2 -44.01 25.3 -43.2 ;
        RECT 24 -44.01 24.1 -43.2 ;
        RECT 22.8 -44.01 22.9 -43.2 ;
        RECT 21.6 -44.01 21.7 -43.2 ;
        RECT 20.4 -44.01 20.5 -43.2 ;
        RECT 19.2 -44.01 19.3 -43.2 ;
        RECT 18 -44.01 18.1 -43.2 ;
        RECT 16.8 -44.01 16.9 -43.2 ;
        RECT 15.6 -44.01 15.7 -43.2 ;
        RECT 14.4 -44.01 14.5 -43.2 ;
        RECT 13.2 -44.01 13.3 -43.2 ;
        RECT 12 -44.01 12.1 -43.2 ;
        RECT 10.8 -44.01 10.9 -43.2 ;
        RECT 9.6 -44.01 9.7 -43.2 ;
        RECT 8.4 -44.01 8.5 -43.2 ;
        RECT 7.2 -44.01 7.3 -43.2 ;
        RECT 6 -44.01 6.1 -43.2 ;
        RECT 4.8 -44.01 4.9 -43.2 ;
        RECT 3.6 -44.01 3.7 -43.2 ;
        RECT 2.4 -44.01 2.5 -43.2 ;
        RECT 1.2 -44.01 1.3 -43.2 ;
        RECT 0 -44.01 0.1 -43.2 ;
        RECT -0.055 -40.435 41.265 -40.315 ;
        RECT 38.4 -40.78 38.5 -39.97 ;
        RECT 37.2 -40.78 37.3 -39.97 ;
        RECT 36 -40.78 36.1 -39.97 ;
        RECT 34.8 -40.78 34.9 -39.97 ;
        RECT 33.6 -40.78 33.7 -39.97 ;
        RECT 32.4 -40.78 32.5 -39.97 ;
        RECT 31.2 -40.78 31.3 -39.97 ;
        RECT 30 -40.78 30.1 -39.97 ;
        RECT 28.8 -40.78 28.9 -39.97 ;
        RECT 27.6 -40.78 27.7 -39.97 ;
        RECT 26.4 -40.78 26.5 -39.97 ;
        RECT 25.2 -40.78 25.3 -39.97 ;
        RECT 24 -40.78 24.1 -39.97 ;
        RECT 22.8 -40.78 22.9 -39.97 ;
        RECT 21.6 -40.78 21.7 -39.97 ;
        RECT 20.4 -40.78 20.5 -39.97 ;
        RECT 19.2 -40.78 19.3 -39.97 ;
        RECT 18 -40.78 18.1 -39.97 ;
        RECT 16.8 -40.78 16.9 -39.97 ;
        RECT 15.6 -40.78 15.7 -39.97 ;
        RECT 14.4 -40.78 14.5 -39.97 ;
        RECT 13.2 -40.78 13.3 -39.97 ;
        RECT 12 -40.78 12.1 -39.97 ;
        RECT 10.8 -40.78 10.9 -39.97 ;
        RECT 9.6 -40.78 9.7 -39.97 ;
        RECT 8.4 -40.78 8.5 -39.97 ;
        RECT 7.2 -40.78 7.3 -39.97 ;
        RECT 6 -40.78 6.1 -39.97 ;
        RECT 4.8 -40.78 4.9 -39.97 ;
        RECT 3.6 -40.78 3.7 -39.97 ;
        RECT 2.4 -40.78 2.5 -39.97 ;
        RECT 1.2 -40.78 1.3 -39.97 ;
        RECT 0 -40.78 0.1 -39.97 ;
        RECT -0.055 -37.205 41.265 -37.085 ;
        RECT 38.4 -37.55 38.5 -36.74 ;
        RECT 37.2 -37.55 37.3 -36.74 ;
        RECT 36 -37.55 36.1 -36.74 ;
        RECT 34.8 -37.55 34.9 -36.74 ;
        RECT 33.6 -37.55 33.7 -36.74 ;
        RECT 32.4 -37.55 32.5 -36.74 ;
        RECT 31.2 -37.55 31.3 -36.74 ;
        RECT 30 -37.55 30.1 -36.74 ;
        RECT 28.8 -37.55 28.9 -36.74 ;
        RECT 27.6 -37.55 27.7 -36.74 ;
        RECT 26.4 -37.55 26.5 -36.74 ;
        RECT 25.2 -37.55 25.3 -36.74 ;
        RECT 24 -37.55 24.1 -36.74 ;
        RECT 22.8 -37.55 22.9 -36.74 ;
        RECT 21.6 -37.55 21.7 -36.74 ;
        RECT 20.4 -37.55 20.5 -36.74 ;
        RECT 19.2 -37.55 19.3 -36.74 ;
        RECT 18 -37.55 18.1 -36.74 ;
        RECT 16.8 -37.55 16.9 -36.74 ;
        RECT 15.6 -37.55 15.7 -36.74 ;
        RECT 14.4 -37.55 14.5 -36.74 ;
        RECT 13.2 -37.55 13.3 -36.74 ;
        RECT 12 -37.55 12.1 -36.74 ;
        RECT 10.8 -37.55 10.9 -36.74 ;
        RECT 9.6 -37.55 9.7 -36.74 ;
        RECT 8.4 -37.55 8.5 -36.74 ;
        RECT 7.2 -37.55 7.3 -36.74 ;
        RECT 6 -37.55 6.1 -36.74 ;
        RECT 4.8 -37.55 4.9 -36.74 ;
        RECT 3.6 -37.55 3.7 -36.74 ;
        RECT 2.4 -37.55 2.5 -36.74 ;
        RECT 1.2 -37.55 1.3 -36.74 ;
        RECT 0 -37.55 0.1 -36.74 ;
        RECT -0.055 -33.975 41.265 -33.855 ;
        RECT 38.4 -34.32 38.5 -33.51 ;
        RECT 37.2 -34.32 37.3 -33.51 ;
        RECT 36 -34.32 36.1 -33.51 ;
        RECT 34.8 -34.32 34.9 -33.51 ;
        RECT 33.6 -34.32 33.7 -33.51 ;
        RECT 32.4 -34.32 32.5 -33.51 ;
        RECT 31.2 -34.32 31.3 -33.51 ;
        RECT 30 -34.32 30.1 -33.51 ;
        RECT 28.8 -34.32 28.9 -33.51 ;
        RECT 27.6 -34.32 27.7 -33.51 ;
        RECT 26.4 -34.32 26.5 -33.51 ;
        RECT 25.2 -34.32 25.3 -33.51 ;
        RECT 24 -34.32 24.1 -33.51 ;
        RECT 22.8 -34.32 22.9 -33.51 ;
        RECT 21.6 -34.32 21.7 -33.51 ;
        RECT 20.4 -34.32 20.5 -33.51 ;
        RECT 19.2 -34.32 19.3 -33.51 ;
        RECT 18 -34.32 18.1 -33.51 ;
        RECT 16.8 -34.32 16.9 -33.51 ;
        RECT 15.6 -34.32 15.7 -33.51 ;
        RECT 14.4 -34.32 14.5 -33.51 ;
        RECT 13.2 -34.32 13.3 -33.51 ;
        RECT 12 -34.32 12.1 -33.51 ;
        RECT 10.8 -34.32 10.9 -33.51 ;
        RECT 9.6 -34.32 9.7 -33.51 ;
        RECT 8.4 -34.32 8.5 -33.51 ;
        RECT 7.2 -34.32 7.3 -33.51 ;
        RECT 6 -34.32 6.1 -33.51 ;
        RECT 4.8 -34.32 4.9 -33.51 ;
        RECT 3.6 -34.32 3.7 -33.51 ;
        RECT 2.4 -34.32 2.5 -33.51 ;
        RECT 1.2 -34.32 1.3 -33.51 ;
        RECT 0 -34.32 0.1 -33.51 ;
        RECT -0.055 -30.745 41.265 -30.625 ;
        RECT 38.4 -31.09 38.5 -30.28 ;
        RECT 37.2 -31.09 37.3 -30.28 ;
        RECT 36 -31.09 36.1 -30.28 ;
        RECT 34.8 -31.09 34.9 -30.28 ;
        RECT 33.6 -31.09 33.7 -30.28 ;
        RECT 32.4 -31.09 32.5 -30.28 ;
        RECT 31.2 -31.09 31.3 -30.28 ;
        RECT 30 -31.09 30.1 -30.28 ;
        RECT 28.8 -31.09 28.9 -30.28 ;
        RECT 27.6 -31.09 27.7 -30.28 ;
        RECT 26.4 -31.09 26.5 -30.28 ;
        RECT 25.2 -31.09 25.3 -30.28 ;
        RECT 24 -31.09 24.1 -30.28 ;
        RECT 22.8 -31.09 22.9 -30.28 ;
        RECT 21.6 -31.09 21.7 -30.28 ;
        RECT 20.4 -31.09 20.5 -30.28 ;
        RECT 19.2 -31.09 19.3 -30.28 ;
        RECT 18 -31.09 18.1 -30.28 ;
        RECT 16.8 -31.09 16.9 -30.28 ;
        RECT 15.6 -31.09 15.7 -30.28 ;
        RECT 14.4 -31.09 14.5 -30.28 ;
        RECT 13.2 -31.09 13.3 -30.28 ;
        RECT 12 -31.09 12.1 -30.28 ;
        RECT 10.8 -31.09 10.9 -30.28 ;
        RECT 9.6 -31.09 9.7 -30.28 ;
        RECT 8.4 -31.09 8.5 -30.28 ;
        RECT 7.2 -31.09 7.3 -30.28 ;
        RECT 6 -31.09 6.1 -30.28 ;
        RECT 4.8 -31.09 4.9 -30.28 ;
        RECT 3.6 -31.09 3.7 -30.28 ;
        RECT 2.4 -31.09 2.5 -30.28 ;
        RECT 1.2 -31.09 1.3 -30.28 ;
        RECT 0 -31.09 0.1 -30.28 ;
        RECT -0.055 -27.515 41.265 -27.395 ;
        RECT 38.4 -27.86 38.5 -27.05 ;
        RECT 37.2 -27.86 37.3 -27.05 ;
        RECT 36 -27.86 36.1 -27.05 ;
        RECT 34.8 -27.86 34.9 -27.05 ;
        RECT 33.6 -27.86 33.7 -27.05 ;
        RECT 32.4 -27.86 32.5 -27.05 ;
        RECT 31.2 -27.86 31.3 -27.05 ;
        RECT 30 -27.86 30.1 -27.05 ;
        RECT 28.8 -27.86 28.9 -27.05 ;
        RECT 27.6 -27.86 27.7 -27.05 ;
        RECT 26.4 -27.86 26.5 -27.05 ;
        RECT 25.2 -27.86 25.3 -27.05 ;
        RECT 24 -27.86 24.1 -27.05 ;
        RECT 22.8 -27.86 22.9 -27.05 ;
        RECT 21.6 -27.86 21.7 -27.05 ;
        RECT 20.4 -27.86 20.5 -27.05 ;
        RECT 19.2 -27.86 19.3 -27.05 ;
        RECT 18 -27.86 18.1 -27.05 ;
        RECT 16.8 -27.86 16.9 -27.05 ;
        RECT 15.6 -27.86 15.7 -27.05 ;
        RECT 14.4 -27.86 14.5 -27.05 ;
        RECT 13.2 -27.86 13.3 -27.05 ;
        RECT 12 -27.86 12.1 -27.05 ;
        RECT 10.8 -27.86 10.9 -27.05 ;
        RECT 9.6 -27.86 9.7 -27.05 ;
        RECT 8.4 -27.86 8.5 -27.05 ;
        RECT 7.2 -27.86 7.3 -27.05 ;
        RECT 6 -27.86 6.1 -27.05 ;
        RECT 4.8 -27.86 4.9 -27.05 ;
        RECT 3.6 -27.86 3.7 -27.05 ;
        RECT 2.4 -27.86 2.5 -27.05 ;
        RECT 1.2 -27.86 1.3 -27.05 ;
        RECT 0 -27.86 0.1 -27.05 ;
        RECT -0.055 -24.285 41.265 -24.165 ;
        RECT 38.4 -24.63 38.5 -23.82 ;
        RECT 37.2 -24.63 37.3 -23.82 ;
        RECT 36 -24.63 36.1 -23.82 ;
        RECT 34.8 -24.63 34.9 -23.82 ;
        RECT 33.6 -24.63 33.7 -23.82 ;
        RECT 32.4 -24.63 32.5 -23.82 ;
        RECT 31.2 -24.63 31.3 -23.82 ;
        RECT 30 -24.63 30.1 -23.82 ;
        RECT 28.8 -24.63 28.9 -23.82 ;
        RECT 27.6 -24.63 27.7 -23.82 ;
        RECT 26.4 -24.63 26.5 -23.82 ;
        RECT 25.2 -24.63 25.3 -23.82 ;
        RECT 24 -24.63 24.1 -23.82 ;
        RECT 22.8 -24.63 22.9 -23.82 ;
        RECT 21.6 -24.63 21.7 -23.82 ;
        RECT 20.4 -24.63 20.5 -23.82 ;
        RECT 19.2 -24.63 19.3 -23.82 ;
        RECT 18 -24.63 18.1 -23.82 ;
        RECT 16.8 -24.63 16.9 -23.82 ;
        RECT 15.6 -24.63 15.7 -23.82 ;
        RECT 14.4 -24.63 14.5 -23.82 ;
        RECT 13.2 -24.63 13.3 -23.82 ;
        RECT 12 -24.63 12.1 -23.82 ;
        RECT 10.8 -24.63 10.9 -23.82 ;
        RECT 9.6 -24.63 9.7 -23.82 ;
        RECT 8.4 -24.63 8.5 -23.82 ;
        RECT 7.2 -24.63 7.3 -23.82 ;
        RECT 6 -24.63 6.1 -23.82 ;
        RECT 4.8 -24.63 4.9 -23.82 ;
        RECT 3.6 -24.63 3.7 -23.82 ;
        RECT 2.4 -24.63 2.5 -23.82 ;
        RECT 1.2 -24.63 1.3 -23.82 ;
        RECT 0 -24.63 0.1 -23.82 ;
        RECT -0.055 -21.055 41.265 -20.935 ;
        RECT 38.4 -21.4 38.5 -20.59 ;
        RECT 37.2 -21.4 37.3 -20.59 ;
        RECT 36 -21.4 36.1 -20.59 ;
        RECT 34.8 -21.4 34.9 -20.59 ;
        RECT 33.6 -21.4 33.7 -20.59 ;
        RECT 32.4 -21.4 32.5 -20.59 ;
        RECT 31.2 -21.4 31.3 -20.59 ;
        RECT 30 -21.4 30.1 -20.59 ;
        RECT 28.8 -21.4 28.9 -20.59 ;
        RECT 27.6 -21.4 27.7 -20.59 ;
        RECT 26.4 -21.4 26.5 -20.59 ;
        RECT 25.2 -21.4 25.3 -20.59 ;
        RECT 24 -21.4 24.1 -20.59 ;
        RECT 22.8 -21.4 22.9 -20.59 ;
        RECT 21.6 -21.4 21.7 -20.59 ;
        RECT 20.4 -21.4 20.5 -20.59 ;
        RECT 19.2 -21.4 19.3 -20.59 ;
        RECT 18 -21.4 18.1 -20.59 ;
        RECT 16.8 -21.4 16.9 -20.59 ;
        RECT 15.6 -21.4 15.7 -20.59 ;
        RECT 14.4 -21.4 14.5 -20.59 ;
        RECT 13.2 -21.4 13.3 -20.59 ;
        RECT 12 -21.4 12.1 -20.59 ;
        RECT 10.8 -21.4 10.9 -20.59 ;
        RECT 9.6 -21.4 9.7 -20.59 ;
        RECT 8.4 -21.4 8.5 -20.59 ;
        RECT 7.2 -21.4 7.3 -20.59 ;
        RECT 6 -21.4 6.1 -20.59 ;
        RECT 4.8 -21.4 4.9 -20.59 ;
        RECT 3.6 -21.4 3.7 -20.59 ;
        RECT 2.4 -21.4 2.5 -20.59 ;
        RECT 1.2 -21.4 1.3 -20.59 ;
        RECT 0 -21.4 0.1 -20.59 ;
        RECT -0.055 -17.825 41.265 -17.705 ;
        RECT 38.4 -18.17 38.5 -17.36 ;
        RECT 37.2 -18.17 37.3 -17.36 ;
        RECT 36 -18.17 36.1 -17.36 ;
        RECT 34.8 -18.17 34.9 -17.36 ;
        RECT 33.6 -18.17 33.7 -17.36 ;
        RECT 32.4 -18.17 32.5 -17.36 ;
        RECT 31.2 -18.17 31.3 -17.36 ;
        RECT 30 -18.17 30.1 -17.36 ;
        RECT 28.8 -18.17 28.9 -17.36 ;
        RECT 27.6 -18.17 27.7 -17.36 ;
        RECT 26.4 -18.17 26.5 -17.36 ;
        RECT 25.2 -18.17 25.3 -17.36 ;
        RECT 24 -18.17 24.1 -17.36 ;
        RECT 22.8 -18.17 22.9 -17.36 ;
        RECT 21.6 -18.17 21.7 -17.36 ;
        RECT 20.4 -18.17 20.5 -17.36 ;
        RECT 19.2 -18.17 19.3 -17.36 ;
        RECT 18 -18.17 18.1 -17.36 ;
        RECT 16.8 -18.17 16.9 -17.36 ;
        RECT 15.6 -18.17 15.7 -17.36 ;
        RECT 14.4 -18.17 14.5 -17.36 ;
        RECT 13.2 -18.17 13.3 -17.36 ;
        RECT 12 -18.17 12.1 -17.36 ;
        RECT 10.8 -18.17 10.9 -17.36 ;
        RECT 9.6 -18.17 9.7 -17.36 ;
        RECT 8.4 -18.17 8.5 -17.36 ;
        RECT 7.2 -18.17 7.3 -17.36 ;
        RECT 6 -18.17 6.1 -17.36 ;
        RECT 4.8 -18.17 4.9 -17.36 ;
        RECT 3.6 -18.17 3.7 -17.36 ;
        RECT 2.4 -18.17 2.5 -17.36 ;
        RECT 1.2 -18.17 1.3 -17.36 ;
        RECT 0 -18.17 0.1 -17.36 ;
        RECT -0.055 -14.595 41.265 -14.475 ;
        RECT 38.4 -14.94 38.5 -14.13 ;
        RECT 37.2 -14.94 37.3 -14.13 ;
        RECT 36 -14.94 36.1 -14.13 ;
        RECT 34.8 -14.94 34.9 -14.13 ;
        RECT 33.6 -14.94 33.7 -14.13 ;
        RECT 32.4 -14.94 32.5 -14.13 ;
        RECT 31.2 -14.94 31.3 -14.13 ;
        RECT 30 -14.94 30.1 -14.13 ;
        RECT 28.8 -14.94 28.9 -14.13 ;
        RECT 27.6 -14.94 27.7 -14.13 ;
        RECT 26.4 -14.94 26.5 -14.13 ;
        RECT 25.2 -14.94 25.3 -14.13 ;
        RECT 24 -14.94 24.1 -14.13 ;
        RECT 22.8 -14.94 22.9 -14.13 ;
        RECT 21.6 -14.94 21.7 -14.13 ;
        RECT 20.4 -14.94 20.5 -14.13 ;
        RECT 19.2 -14.94 19.3 -14.13 ;
        RECT 18 -14.94 18.1 -14.13 ;
        RECT 16.8 -14.94 16.9 -14.13 ;
        RECT 15.6 -14.94 15.7 -14.13 ;
        RECT 14.4 -14.94 14.5 -14.13 ;
        RECT 13.2 -14.94 13.3 -14.13 ;
        RECT 12 -14.94 12.1 -14.13 ;
        RECT 10.8 -14.94 10.9 -14.13 ;
        RECT 9.6 -14.94 9.7 -14.13 ;
        RECT 8.4 -14.94 8.5 -14.13 ;
        RECT 7.2 -14.94 7.3 -14.13 ;
        RECT 6 -14.94 6.1 -14.13 ;
        RECT 4.8 -14.94 4.9 -14.13 ;
        RECT 3.6 -14.94 3.7 -14.13 ;
        RECT 2.4 -14.94 2.5 -14.13 ;
        RECT 1.2 -14.94 1.3 -14.13 ;
        RECT 0 -14.94 0.1 -14.13 ;
        RECT -0.055 -11.365 41.265 -11.245 ;
        RECT 38.4 -11.71 38.5 -10.9 ;
        RECT 37.2 -11.71 37.3 -10.9 ;
        RECT 36 -11.71 36.1 -10.9 ;
        RECT 34.8 -11.71 34.9 -10.9 ;
        RECT 33.6 -11.71 33.7 -10.9 ;
        RECT 32.4 -11.71 32.5 -10.9 ;
        RECT 31.2 -11.71 31.3 -10.9 ;
        RECT 30 -11.71 30.1 -10.9 ;
        RECT 28.8 -11.71 28.9 -10.9 ;
        RECT 27.6 -11.71 27.7 -10.9 ;
        RECT 26.4 -11.71 26.5 -10.9 ;
        RECT 25.2 -11.71 25.3 -10.9 ;
        RECT 24 -11.71 24.1 -10.9 ;
        RECT 22.8 -11.71 22.9 -10.9 ;
        RECT 21.6 -11.71 21.7 -10.9 ;
        RECT 20.4 -11.71 20.5 -10.9 ;
        RECT 19.2 -11.71 19.3 -10.9 ;
        RECT 18 -11.71 18.1 -10.9 ;
        RECT 16.8 -11.71 16.9 -10.9 ;
        RECT 15.6 -11.71 15.7 -10.9 ;
        RECT 14.4 -11.71 14.5 -10.9 ;
        RECT 13.2 -11.71 13.3 -10.9 ;
        RECT 12 -11.71 12.1 -10.9 ;
        RECT 10.8 -11.71 10.9 -10.9 ;
        RECT 9.6 -11.71 9.7 -10.9 ;
        RECT 8.4 -11.71 8.5 -10.9 ;
        RECT 7.2 -11.71 7.3 -10.9 ;
        RECT 6 -11.71 6.1 -10.9 ;
        RECT 4.8 -11.71 4.9 -10.9 ;
        RECT 3.6 -11.71 3.7 -10.9 ;
        RECT 2.4 -11.71 2.5 -10.9 ;
        RECT 1.2 -11.71 1.3 -10.9 ;
        RECT 0 -11.71 0.1 -10.9 ;
        RECT -0.055 -8.135 41.265 -8.015 ;
        RECT 38.4 -8.48 38.5 -7.67 ;
        RECT 37.2 -8.48 37.3 -7.67 ;
        RECT 36 -8.48 36.1 -7.67 ;
        RECT 34.8 -8.48 34.9 -7.67 ;
        RECT 33.6 -8.48 33.7 -7.67 ;
        RECT 32.4 -8.48 32.5 -7.67 ;
        RECT 31.2 -8.48 31.3 -7.67 ;
        RECT 30 -8.48 30.1 -7.67 ;
        RECT 28.8 -8.48 28.9 -7.67 ;
        RECT 27.6 -8.48 27.7 -7.67 ;
        RECT 26.4 -8.48 26.5 -7.67 ;
        RECT 25.2 -8.48 25.3 -7.67 ;
        RECT 24 -8.48 24.1 -7.67 ;
        RECT 22.8 -8.48 22.9 -7.67 ;
        RECT 21.6 -8.48 21.7 -7.67 ;
        RECT 20.4 -8.48 20.5 -7.67 ;
        RECT 19.2 -8.48 19.3 -7.67 ;
        RECT 18 -8.48 18.1 -7.67 ;
        RECT 16.8 -8.48 16.9 -7.67 ;
        RECT 15.6 -8.48 15.7 -7.67 ;
        RECT 14.4 -8.48 14.5 -7.67 ;
        RECT 13.2 -8.48 13.3 -7.67 ;
        RECT 12 -8.48 12.1 -7.67 ;
        RECT 10.8 -8.48 10.9 -7.67 ;
        RECT 9.6 -8.48 9.7 -7.67 ;
        RECT 8.4 -8.48 8.5 -7.67 ;
        RECT 7.2 -8.48 7.3 -7.67 ;
        RECT 6 -8.48 6.1 -7.67 ;
        RECT 4.8 -8.48 4.9 -7.67 ;
        RECT 3.6 -8.48 3.7 -7.67 ;
        RECT 2.4 -8.48 2.5 -7.67 ;
        RECT 1.2 -8.48 1.3 -7.67 ;
        RECT 0 -8.48 0.1 -7.67 ;
        RECT -0.055 -4.905 41.265 -4.785 ;
        RECT 38.4 -5.25 38.5 -4.44 ;
        RECT 37.2 -5.25 37.3 -4.44 ;
        RECT 36 -5.25 36.1 -4.44 ;
        RECT 34.8 -5.25 34.9 -4.44 ;
        RECT 33.6 -5.25 33.7 -4.44 ;
        RECT 32.4 -5.25 32.5 -4.44 ;
        RECT 31.2 -5.25 31.3 -4.44 ;
        RECT 30 -5.25 30.1 -4.44 ;
        RECT 28.8 -5.25 28.9 -4.44 ;
        RECT 27.6 -5.25 27.7 -4.44 ;
        RECT 26.4 -5.25 26.5 -4.44 ;
        RECT 25.2 -5.25 25.3 -4.44 ;
        RECT 24 -5.25 24.1 -4.44 ;
        RECT 22.8 -5.25 22.9 -4.44 ;
        RECT 21.6 -5.25 21.7 -4.44 ;
        RECT 20.4 -5.25 20.5 -4.44 ;
        RECT 19.2 -5.25 19.3 -4.44 ;
        RECT 18 -5.25 18.1 -4.44 ;
        RECT 16.8 -5.25 16.9 -4.44 ;
        RECT 15.6 -5.25 15.7 -4.44 ;
        RECT 14.4 -5.25 14.5 -4.44 ;
        RECT 13.2 -5.25 13.3 -4.44 ;
        RECT 12 -5.25 12.1 -4.44 ;
        RECT 10.8 -5.25 10.9 -4.44 ;
        RECT 9.6 -5.25 9.7 -4.44 ;
        RECT 8.4 -5.25 8.5 -4.44 ;
        RECT 7.2 -5.25 7.3 -4.44 ;
        RECT 6 -5.25 6.1 -4.44 ;
        RECT 4.8 -5.25 4.9 -4.44 ;
        RECT 3.6 -5.25 3.7 -4.44 ;
        RECT 2.4 -5.25 2.5 -4.44 ;
        RECT 1.2 -5.25 1.3 -4.44 ;
        RECT 0 -5.25 0.1 -4.44 ;
        RECT -0.055 -1.675 41.265 -1.555 ;
        RECT 38.4 -2.02 38.5 -1.21 ;
        RECT 37.2 -2.02 37.3 -1.21 ;
        RECT 36 -2.02 36.1 -1.21 ;
        RECT 34.8 -2.02 34.9 -1.21 ;
        RECT 33.6 -2.02 33.7 -1.21 ;
        RECT 32.4 -2.02 32.5 -1.21 ;
        RECT 31.2 -2.02 31.3 -1.21 ;
        RECT 30 -2.02 30.1 -1.21 ;
        RECT 28.8 -2.02 28.9 -1.21 ;
        RECT 27.6 -2.02 27.7 -1.21 ;
        RECT 26.4 -2.02 26.5 -1.21 ;
        RECT 25.2 -2.02 25.3 -1.21 ;
        RECT 24 -2.02 24.1 -1.21 ;
        RECT 22.8 -2.02 22.9 -1.21 ;
        RECT 21.6 -2.02 21.7 -1.21 ;
        RECT 20.4 -2.02 20.5 -1.21 ;
        RECT 19.2 -2.02 19.3 -1.21 ;
        RECT 18 -2.02 18.1 -1.21 ;
        RECT 16.8 -2.02 16.9 -1.21 ;
        RECT 15.6 -2.02 15.7 -1.21 ;
        RECT 14.4 -2.02 14.5 -1.21 ;
        RECT 13.2 -2.02 13.3 -1.21 ;
        RECT 12 -2.02 12.1 -1.21 ;
        RECT 10.8 -2.02 10.9 -1.21 ;
        RECT 9.6 -2.02 9.7 -1.21 ;
        RECT 8.4 -2.02 8.5 -1.21 ;
        RECT 7.2 -2.02 7.3 -1.21 ;
        RECT 6 -2.02 6.1 -1.21 ;
        RECT 4.8 -2.02 4.9 -1.21 ;
        RECT 3.6 -2.02 3.7 -1.21 ;
        RECT 2.4 -2.02 2.5 -1.21 ;
        RECT 1.2 -2.02 1.3 -1.21 ;
        RECT 0 -2.02 0.1 -1.21 ;
        RECT -0.055 1.555 41.265 1.675 ;
        RECT 38.4 1.21 38.5 1.675 ;
        RECT 37.2 1.21 37.3 1.675 ;
        RECT 36 1.21 36.1 1.675 ;
        RECT 34.8 1.21 34.9 1.675 ;
        RECT 33.6 1.21 33.7 1.675 ;
        RECT 32.4 1.21 32.5 1.675 ;
        RECT 31.2 1.21 31.3 1.675 ;
        RECT 30 1.21 30.1 1.675 ;
        RECT 28.8 1.21 28.9 1.675 ;
        RECT 27.6 1.21 27.7 1.675 ;
        RECT 26.4 1.21 26.5 1.675 ;
        RECT 25.2 1.21 25.3 1.675 ;
        RECT 24 1.21 24.1 1.675 ;
        RECT 22.8 1.21 22.9 1.675 ;
        RECT 21.6 1.21 21.7 1.675 ;
        RECT 20.4 1.21 20.5 1.675 ;
        RECT 19.2 1.21 19.3 1.675 ;
        RECT 18 1.21 18.1 1.675 ;
        RECT 16.8 1.21 16.9 1.675 ;
        RECT 15.6 1.21 15.7 1.675 ;
        RECT 14.4 1.21 14.5 1.675 ;
        RECT 13.2 1.21 13.3 1.675 ;
        RECT 12 1.21 12.1 1.675 ;
        RECT 10.8 1.21 10.9 1.675 ;
        RECT 9.6 1.21 9.7 1.675 ;
        RECT 8.4 1.21 8.5 1.675 ;
        RECT 7.2 1.21 7.3 1.675 ;
        RECT 6 1.21 6.1 1.675 ;
        RECT 4.8 1.21 4.9 1.675 ;
        RECT 3.6 1.21 3.7 1.675 ;
        RECT 2.4 1.21 2.5 1.675 ;
        RECT 1.2 1.21 1.3 1.675 ;
        RECT 0 1.21 0.1 1.675 ;
        RECT 0.04 3.42 41.265 3.8 ;
        RECT 38.275 2.175 38.375 3.8 ;
        RECT 37.325 2.175 37.425 3.8 ;
        RECT 37.075 2.175 37.175 3.8 ;
        RECT 36.125 2.175 36.225 3.8 ;
        RECT 35.875 2.175 35.975 3.8 ;
        RECT 34.925 2.175 35.025 3.8 ;
        RECT 34.675 2.175 34.775 3.8 ;
        RECT 33.725 2.175 33.825 3.8 ;
        RECT 33.475 2.175 33.575 3.8 ;
        RECT 32.525 2.175 32.625 3.8 ;
        RECT 32.275 2.175 32.375 3.8 ;
        RECT 31.325 2.175 31.425 3.8 ;
        RECT 31.075 2.175 31.175 3.8 ;
        RECT 30.125 2.175 30.225 3.8 ;
        RECT 29.875 2.175 29.975 3.8 ;
        RECT 28.925 2.175 29.025 3.8 ;
        RECT 28.675 2.175 28.775 3.8 ;
        RECT 27.725 2.175 27.825 3.8 ;
        RECT 27.475 2.175 27.575 3.8 ;
        RECT 26.525 2.175 26.625 3.8 ;
        RECT 26.275 2.175 26.375 3.8 ;
        RECT 25.325 2.175 25.425 3.8 ;
        RECT 25.075 2.175 25.175 3.8 ;
        RECT 24.125 2.175 24.225 3.8 ;
        RECT 23.875 2.175 23.975 3.8 ;
        RECT 22.925 2.175 23.025 3.8 ;
        RECT 22.675 2.175 22.775 3.8 ;
        RECT 21.725 2.175 21.825 3.8 ;
        RECT 21.475 2.175 21.575 3.8 ;
        RECT 20.525 2.175 20.625 3.8 ;
        RECT 20.275 2.175 20.375 3.8 ;
        RECT 19.325 2.175 19.425 3.8 ;
        RECT 19.075 2.175 19.175 3.8 ;
        RECT 18.125 2.175 18.225 3.8 ;
        RECT 17.875 2.175 17.975 3.8 ;
        RECT 16.925 2.175 17.025 3.8 ;
        RECT 16.675 2.175 16.775 3.8 ;
        RECT 15.725 2.175 15.825 3.8 ;
        RECT 15.475 2.175 15.575 3.8 ;
        RECT 14.525 2.175 14.625 3.8 ;
        RECT 14.275 2.175 14.375 3.8 ;
        RECT 13.325 2.175 13.425 3.8 ;
        RECT 13.075 2.175 13.175 3.8 ;
        RECT 12.125 2.175 12.225 3.8 ;
        RECT 11.875 2.175 11.975 3.8 ;
        RECT 10.925 2.175 11.025 3.8 ;
        RECT 10.675 2.175 10.775 3.8 ;
        RECT 9.725 2.175 9.825 3.8 ;
        RECT 9.475 2.175 9.575 3.8 ;
        RECT 8.525 2.175 8.625 3.8 ;
        RECT 8.275 2.175 8.375 3.8 ;
        RECT 7.325 2.175 7.425 3.8 ;
        RECT 7.075 2.175 7.175 3.8 ;
        RECT 6.125 2.175 6.225 3.8 ;
        RECT 5.875 2.175 5.975 3.8 ;
        RECT 4.925 2.175 5.025 3.8 ;
        RECT 4.675 2.175 4.775 3.8 ;
        RECT 3.725 2.175 3.825 3.8 ;
        RECT 3.475 2.175 3.575 3.8 ;
        RECT 2.525 2.175 2.625 3.8 ;
        RECT 2.275 2.175 2.375 3.8 ;
        RECT 1.325 2.175 1.425 3.8 ;
        RECT 1.075 2.175 1.175 3.8 ;
        RECT 0.125 2.175 0.225 3.8 ;
        RECT -31.525 -50.405 -0.585 -49.725 ;
        RECT -1.025 -51.215 -0.925 -48.915 ;
        RECT -1.545 -51.215 -1.445 -48.915 ;
        RECT -2.325 -51.215 -2.225 -48.915 ;
        RECT -2.845 -51.215 -2.745 -48.915 ;
        RECT -3.625 -51.215 -3.525 -48.915 ;
        RECT -4.145 -51.215 -4.045 -48.915 ;
        RECT -4.925 -51.215 -4.825 -48.915 ;
        RECT -5.445 -51.215 -5.345 -48.915 ;
        RECT -6.225 -51.215 -6.125 -48.915 ;
        RECT -6.745 -51.215 -6.645 -48.915 ;
        RECT -7.525 -51.215 -7.425 -48.915 ;
        RECT -8.045 -51.215 -7.945 -48.915 ;
        RECT -8.825 -51.215 -8.725 -48.915 ;
        RECT -9.345 -51.215 -9.245 -48.915 ;
        RECT -10.125 -51.215 -10.025 -48.915 ;
        RECT -10.645 -51.215 -10.545 -48.915 ;
        RECT -11.425 -50.405 -11.325 -48.915 ;
        RECT -11.945 -50.405 -11.845 -48.915 ;
        RECT -12.725 -50.405 -12.625 -48.915 ;
        RECT -13.245 -50.405 -13.145 -48.915 ;
        RECT -14.025 -50.405 -13.925 -48.915 ;
        RECT -14.545 -50.405 -14.445 -48.915 ;
        RECT -15.325 -50.405 -15.225 -48.915 ;
        RECT -15.845 -50.405 -15.745 -48.915 ;
        RECT -16.625 -50.405 -16.525 -48.915 ;
        RECT -17.145 -50.405 -17.045 -48.915 ;
        RECT -17.925 -50.405 -17.825 -48.915 ;
        RECT -18.445 -50.405 -18.345 -48.915 ;
        RECT -19.225 -50.405 -19.125 -48.915 ;
        RECT -19.745 -50.405 -19.645 -48.915 ;
        RECT -20.525 -50.405 -20.425 -48.915 ;
        RECT -21.045 -50.405 -20.945 -48.915 ;
        RECT -21.825 -50.405 -21.725 -48.915 ;
        RECT -22.345 -50.405 -22.245 -48.915 ;
        RECT -23.125 -50.405 -23.025 -48.915 ;
        RECT -23.645 -50.405 -23.545 -48.915 ;
        RECT -24.425 -50.405 -24.325 -48.915 ;
        RECT -24.945 -50.405 -24.845 -48.915 ;
        RECT -25.725 -50.405 -25.625 -48.915 ;
        RECT -26.245 -50.405 -26.145 -48.915 ;
        RECT -31.525 -37.485 -0.585 -36.805 ;
        RECT -1.025 -38.295 -0.925 -35.995 ;
        RECT -1.545 -38.295 -1.445 -35.995 ;
        RECT -2.325 -38.295 -2.225 -35.995 ;
        RECT -2.845 -38.295 -2.745 -35.995 ;
        RECT -3.625 -38.295 -3.525 -35.995 ;
        RECT -4.145 -38.295 -4.045 -35.995 ;
        RECT -4.925 -38.295 -4.825 -35.995 ;
        RECT -5.445 -38.295 -5.345 -35.995 ;
        RECT -6.225 -38.295 -6.125 -35.995 ;
        RECT -6.745 -38.295 -6.645 -35.995 ;
        RECT -7.525 -38.295 -7.425 -35.995 ;
        RECT -8.045 -38.295 -7.945 -35.995 ;
        RECT -8.825 -38.295 -8.725 -35.995 ;
        RECT -9.345 -38.295 -9.245 -35.995 ;
        RECT -10.125 -38.295 -10.025 -35.995 ;
        RECT -10.645 -38.295 -10.545 -35.995 ;
        RECT -11.425 -38.295 -11.325 -35.995 ;
        RECT -11.945 -38.295 -11.845 -35.995 ;
        RECT -12.725 -38.295 -12.625 -35.995 ;
        RECT -13.245 -38.295 -13.145 -35.995 ;
        RECT -14.025 -38.295 -13.925 -35.995 ;
        RECT -14.545 -38.295 -14.445 -35.995 ;
        RECT -15.325 -38.295 -15.225 -35.995 ;
        RECT -15.845 -38.295 -15.745 -35.995 ;
        RECT -16.625 -38.295 -16.525 -35.995 ;
        RECT -17.145 -38.295 -17.045 -35.995 ;
        RECT -17.925 -38.295 -17.825 -35.995 ;
        RECT -18.445 -38.295 -18.345 -35.995 ;
        RECT -19.225 -38.295 -19.125 -35.995 ;
        RECT -19.745 -38.295 -19.645 -35.995 ;
        RECT -20.525 -38.295 -20.425 -35.995 ;
        RECT -21.045 -38.295 -20.945 -35.995 ;
        RECT -21.825 -38.295 -21.725 -35.995 ;
        RECT -22.345 -38.295 -22.245 -35.995 ;
        RECT -23.125 -38.295 -23.025 -35.995 ;
        RECT -23.645 -38.295 -23.545 -35.995 ;
        RECT -24.425 -38.295 -24.325 -35.995 ;
        RECT -24.945 -38.295 -24.845 -35.995 ;
        RECT -25.725 -38.295 -25.625 -35.995 ;
        RECT -26.245 -38.295 -26.145 -35.995 ;
        RECT -31.525 -24.565 -0.585 -23.885 ;
        RECT -1.025 -25.375 -0.925 -23.075 ;
        RECT -1.545 -25.375 -1.445 -23.075 ;
        RECT -2.325 -25.375 -2.225 -23.075 ;
        RECT -2.845 -25.375 -2.745 -23.075 ;
        RECT -3.625 -25.375 -3.525 -23.075 ;
        RECT -4.145 -25.375 -4.045 -23.075 ;
        RECT -4.925 -25.375 -4.825 -23.075 ;
        RECT -5.445 -25.375 -5.345 -23.075 ;
        RECT -6.225 -25.375 -6.125 -23.075 ;
        RECT -6.745 -25.375 -6.645 -23.075 ;
        RECT -7.525 -25.375 -7.425 -23.075 ;
        RECT -8.045 -25.375 -7.945 -23.075 ;
        RECT -8.825 -25.375 -8.725 -23.075 ;
        RECT -9.345 -25.375 -9.245 -23.075 ;
        RECT -10.125 -25.375 -10.025 -23.075 ;
        RECT -10.645 -25.375 -10.545 -23.075 ;
        RECT -11.425 -25.375 -11.325 -23.075 ;
        RECT -11.945 -25.375 -11.845 -23.075 ;
        RECT -12.725 -25.375 -12.625 -23.075 ;
        RECT -13.245 -25.375 -13.145 -23.075 ;
        RECT -14.025 -25.375 -13.925 -23.075 ;
        RECT -14.545 -25.375 -14.445 -23.075 ;
        RECT -15.325 -25.375 -15.225 -23.075 ;
        RECT -15.845 -25.375 -15.745 -23.075 ;
        RECT -16.625 -25.375 -16.525 -23.075 ;
        RECT -17.145 -25.375 -17.045 -23.075 ;
        RECT -17.925 -25.375 -17.825 -23.075 ;
        RECT -18.445 -25.375 -18.345 -23.075 ;
        RECT -19.225 -25.375 -19.125 -23.075 ;
        RECT -19.745 -25.375 -19.645 -23.075 ;
        RECT -20.525 -25.375 -20.425 -23.075 ;
        RECT -21.045 -25.375 -20.945 -23.075 ;
        RECT -21.825 -25.375 -21.725 -23.075 ;
        RECT -22.345 -25.375 -22.245 -23.075 ;
        RECT -23.125 -25.375 -23.025 -23.075 ;
        RECT -23.645 -25.375 -23.545 -23.075 ;
        RECT -24.425 -25.375 -24.325 -23.075 ;
        RECT -24.945 -25.375 -24.845 -23.075 ;
        RECT -25.725 -25.375 -25.625 -23.075 ;
        RECT -26.245 -25.375 -26.145 -23.075 ;
        RECT -31.525 -11.645 -0.585 -10.965 ;
        RECT -1.025 -12.455 -0.925 -10.155 ;
        RECT -1.545 -12.455 -1.445 -10.155 ;
        RECT -2.325 -12.455 -2.225 -10.155 ;
        RECT -2.845 -12.455 -2.745 -10.155 ;
        RECT -3.625 -12.455 -3.525 -10.155 ;
        RECT -4.145 -12.455 -4.045 -10.155 ;
        RECT -4.925 -12.455 -4.825 -10.155 ;
        RECT -5.445 -12.455 -5.345 -10.155 ;
        RECT -6.225 -12.455 -6.125 -10.155 ;
        RECT -6.745 -12.455 -6.645 -10.155 ;
        RECT -7.525 -12.455 -7.425 -10.155 ;
        RECT -8.045 -12.455 -7.945 -10.155 ;
        RECT -8.825 -12.455 -8.725 -10.155 ;
        RECT -9.345 -12.455 -9.245 -10.155 ;
        RECT -10.125 -12.455 -10.025 -10.155 ;
        RECT -10.645 -12.455 -10.545 -10.155 ;
        RECT -11.425 -12.455 -11.325 -10.155 ;
        RECT -11.945 -12.455 -11.845 -10.155 ;
        RECT -12.725 -12.455 -12.625 -10.155 ;
        RECT -13.245 -12.455 -13.145 -10.155 ;
        RECT -14.025 -12.455 -13.925 -10.155 ;
        RECT -14.545 -12.455 -14.445 -10.155 ;
        RECT -15.325 -12.455 -15.225 -10.155 ;
        RECT -15.845 -12.455 -15.745 -10.155 ;
        RECT -16.625 -12.455 -16.525 -10.155 ;
        RECT -17.145 -12.455 -17.045 -10.155 ;
        RECT -17.925 -12.455 -17.825 -10.155 ;
        RECT -18.445 -12.455 -18.345 -10.155 ;
        RECT -19.225 -12.455 -19.125 -10.155 ;
        RECT -19.745 -12.455 -19.645 -10.155 ;
        RECT -20.525 -12.455 -20.425 -10.155 ;
        RECT -21.045 -12.455 -20.945 -10.155 ;
        RECT -21.825 -12.455 -21.725 -10.155 ;
        RECT -22.345 -12.455 -22.245 -10.155 ;
        RECT -23.125 -12.455 -23.025 -10.155 ;
        RECT -23.645 -12.455 -23.545 -10.155 ;
        RECT -24.425 -12.455 -24.325 -10.155 ;
        RECT -24.945 -12.455 -24.845 -10.155 ;
        RECT -25.725 -12.455 -25.625 -10.155 ;
        RECT -26.245 -12.455 -26.145 -10.155 ;
        RECT -31.525 1.275 -0.585 1.955 ;
        RECT -1.025 0.465 -0.925 1.955 ;
        RECT -1.545 0.465 -1.445 1.955 ;
        RECT -2.325 0.465 -2.225 1.955 ;
        RECT -2.845 0.465 -2.745 1.955 ;
        RECT -3.625 0.465 -3.525 1.955 ;
        RECT -4.145 0.465 -4.045 1.955 ;
        RECT -4.925 0.465 -4.825 1.955 ;
        RECT -5.445 0.465 -5.345 1.955 ;
        RECT -5.885 1.275 -5.785 2.59 ;
        RECT -6.225 0.465 -6.125 1.955 ;
        RECT -6.445 1.275 -6.345 2.59 ;
        RECT -6.745 0.465 -6.645 1.955 ;
        RECT -7.525 0.465 -7.425 1.955 ;
        RECT -8.045 0.465 -7.945 1.955 ;
        RECT -8.825 0.465 -8.725 1.955 ;
        RECT -9.345 0.465 -9.245 1.955 ;
        RECT -10.125 0.465 -10.025 1.955 ;
        RECT -10.645 0.465 -10.545 1.955 ;
        RECT -11.425 0.465 -11.325 1.955 ;
        RECT -11.945 0.465 -11.845 1.955 ;
        RECT -12.725 0.465 -12.625 1.955 ;
        RECT -13.245 0.465 -13.145 1.955 ;
        RECT -14.025 0.465 -13.925 1.955 ;
        RECT -14.545 0.465 -14.445 1.955 ;
        RECT -15.325 0.465 -15.225 1.955 ;
        RECT -15.845 0.465 -15.745 1.955 ;
        RECT -16.625 0.465 -16.525 1.955 ;
        RECT -17.145 0.465 -17.045 1.955 ;
        RECT -17.925 0.465 -17.825 1.955 ;
        RECT -18.445 0.465 -18.345 1.955 ;
        RECT -19.225 0.465 -19.125 1.955 ;
        RECT -19.745 0.465 -19.645 1.955 ;
        RECT -20.525 0.465 -20.425 1.955 ;
        RECT -21.045 0.465 -20.945 1.955 ;
        RECT -21.825 0.465 -21.725 1.955 ;
        RECT -22.345 0.465 -22.245 1.955 ;
        RECT -23.125 0.465 -23.025 1.955 ;
        RECT -23.645 0.465 -23.545 1.955 ;
        RECT -24.425 0.465 -24.325 1.955 ;
        RECT -24.945 0.465 -24.845 1.955 ;
        RECT -25.725 0.465 -25.625 1.955 ;
        RECT -26.245 0.465 -26.145 1.955 ;
        RECT -27.125 1.275 -27.025 2.645 ;
        RECT -27.725 1.275 -27.625 2.645 ;
        RECT -28.325 1.275 -28.225 2.645 ;
        RECT -28.925 1.275 -28.825 2.645 ;
        RECT -29.525 1.275 -29.425 2.645 ;
        RECT -31.525 -59.845 -10.965 -59.165 ;
        RECT -11.525 -59.845 -11.425 -58.475 ;
        RECT -12.125 -59.845 -12.025 -58.475 ;
      LAYER V1 ;
        RECT -31.42 1.795 -31.32 1.895 ;
        RECT -31.42 1.565 -31.32 1.665 ;
        RECT -31.42 1.335 -31.32 1.435 ;
        RECT -31.42 -11.125 -31.32 -11.025 ;
        RECT -31.42 -11.355 -31.32 -11.255 ;
        RECT -31.42 -11.585 -31.32 -11.485 ;
        RECT -31.42 -24.045 -31.32 -23.945 ;
        RECT -31.42 -24.275 -31.32 -24.175 ;
        RECT -31.42 -24.505 -31.32 -24.405 ;
        RECT -31.42 -36.965 -31.32 -36.865 ;
        RECT -31.42 -37.195 -31.32 -37.095 ;
        RECT -31.42 -37.425 -31.32 -37.325 ;
        RECT -31.42 -49.885 -31.32 -49.785 ;
        RECT -31.42 -50.115 -31.32 -50.015 ;
        RECT -31.42 -50.345 -31.32 -50.245 ;
        RECT -31.42 -59.325 -31.32 -59.225 ;
        RECT -31.42 -59.555 -31.32 -59.455 ;
        RECT -31.42 -59.785 -31.32 -59.685 ;
        RECT -31.42 -66.11 -31.32 -66.01 ;
        RECT -31.42 -66.34 -31.32 -66.24 ;
        RECT -31.42 -66.57 -31.32 -66.47 ;
        RECT -31.42 -66.8 -31.32 -66.7 ;
        RECT -31.42 -67.03 -31.32 -66.93 ;
        RECT -31.42 -67.26 -31.32 -67.16 ;
        RECT -31.42 -67.49 -31.32 -67.39 ;
        RECT -31.42 -67.72 -31.32 -67.62 ;
        RECT -31.42 -67.95 -31.32 -67.85 ;
        RECT -31.42 -68.18 -31.32 -68.08 ;
        RECT -31.42 -68.41 -31.32 -68.31 ;
        RECT -31.42 -68.64 -31.32 -68.54 ;
        RECT -31.19 1.795 -31.09 1.895 ;
        RECT -31.19 1.565 -31.09 1.665 ;
        RECT -31.19 1.335 -31.09 1.435 ;
        RECT -31.19 -11.125 -31.09 -11.025 ;
        RECT -31.19 -11.355 -31.09 -11.255 ;
        RECT -31.19 -11.585 -31.09 -11.485 ;
        RECT -31.19 -24.045 -31.09 -23.945 ;
        RECT -31.19 -24.275 -31.09 -24.175 ;
        RECT -31.19 -24.505 -31.09 -24.405 ;
        RECT -31.19 -36.965 -31.09 -36.865 ;
        RECT -31.19 -37.195 -31.09 -37.095 ;
        RECT -31.19 -37.425 -31.09 -37.325 ;
        RECT -31.19 -49.885 -31.09 -49.785 ;
        RECT -31.19 -50.115 -31.09 -50.015 ;
        RECT -31.19 -50.345 -31.09 -50.245 ;
        RECT -31.19 -59.325 -31.09 -59.225 ;
        RECT -31.19 -59.555 -31.09 -59.455 ;
        RECT -31.19 -59.785 -31.09 -59.685 ;
        RECT -31.19 -66.11 -31.09 -66.01 ;
        RECT -31.19 -66.34 -31.09 -66.24 ;
        RECT -31.19 -66.57 -31.09 -66.47 ;
        RECT -31.19 -66.8 -31.09 -66.7 ;
        RECT -31.19 -67.03 -31.09 -66.93 ;
        RECT -31.19 -67.26 -31.09 -67.16 ;
        RECT -31.19 -67.49 -31.09 -67.39 ;
        RECT -31.19 -67.72 -31.09 -67.62 ;
        RECT -31.19 -67.95 -31.09 -67.85 ;
        RECT -31.19 -68.18 -31.09 -68.08 ;
        RECT -31.19 -68.41 -31.09 -68.31 ;
        RECT -31.19 -68.64 -31.09 -68.54 ;
        RECT -30.96 1.795 -30.86 1.895 ;
        RECT -30.96 1.565 -30.86 1.665 ;
        RECT -30.96 1.335 -30.86 1.435 ;
        RECT -30.96 -11.125 -30.86 -11.025 ;
        RECT -30.96 -11.355 -30.86 -11.255 ;
        RECT -30.96 -11.585 -30.86 -11.485 ;
        RECT -30.96 -24.045 -30.86 -23.945 ;
        RECT -30.96 -24.275 -30.86 -24.175 ;
        RECT -30.96 -24.505 -30.86 -24.405 ;
        RECT -30.96 -36.965 -30.86 -36.865 ;
        RECT -30.96 -37.195 -30.86 -37.095 ;
        RECT -30.96 -37.425 -30.86 -37.325 ;
        RECT -30.96 -49.885 -30.86 -49.785 ;
        RECT -30.96 -50.115 -30.86 -50.015 ;
        RECT -30.96 -50.345 -30.86 -50.245 ;
        RECT -30.96 -59.325 -30.86 -59.225 ;
        RECT -30.96 -59.555 -30.86 -59.455 ;
        RECT -30.96 -59.785 -30.86 -59.685 ;
        RECT -30.96 -66.11 -30.86 -66.01 ;
        RECT -30.96 -66.34 -30.86 -66.24 ;
        RECT -30.96 -66.57 -30.86 -66.47 ;
        RECT -30.96 -66.8 -30.86 -66.7 ;
        RECT -30.96 -67.03 -30.86 -66.93 ;
        RECT -30.96 -67.26 -30.86 -67.16 ;
        RECT -30.96 -67.49 -30.86 -67.39 ;
        RECT -30.96 -67.72 -30.86 -67.62 ;
        RECT -30.96 -67.95 -30.86 -67.85 ;
        RECT -30.96 -68.18 -30.86 -68.08 ;
        RECT -30.96 -68.41 -30.86 -68.31 ;
        RECT -30.96 -68.64 -30.86 -68.54 ;
        RECT -30.73 1.795 -30.63 1.895 ;
        RECT -30.73 1.565 -30.63 1.665 ;
        RECT -30.73 1.335 -30.63 1.435 ;
        RECT -30.73 -11.125 -30.63 -11.025 ;
        RECT -30.73 -11.355 -30.63 -11.255 ;
        RECT -30.73 -11.585 -30.63 -11.485 ;
        RECT -30.73 -24.045 -30.63 -23.945 ;
        RECT -30.73 -24.275 -30.63 -24.175 ;
        RECT -30.73 -24.505 -30.63 -24.405 ;
        RECT -30.73 -36.965 -30.63 -36.865 ;
        RECT -30.73 -37.195 -30.63 -37.095 ;
        RECT -30.73 -37.425 -30.63 -37.325 ;
        RECT -30.73 -49.885 -30.63 -49.785 ;
        RECT -30.73 -50.115 -30.63 -50.015 ;
        RECT -30.73 -50.345 -30.63 -50.245 ;
        RECT -30.73 -59.325 -30.63 -59.225 ;
        RECT -30.73 -59.555 -30.63 -59.455 ;
        RECT -30.73 -59.785 -30.63 -59.685 ;
        RECT -30.73 -66.11 -30.63 -66.01 ;
        RECT -30.73 -66.34 -30.63 -66.24 ;
        RECT -30.73 -66.57 -30.63 -66.47 ;
        RECT -30.73 -66.8 -30.63 -66.7 ;
        RECT -30.73 -67.03 -30.63 -66.93 ;
        RECT -30.73 -67.26 -30.63 -67.16 ;
        RECT -30.73 -67.49 -30.63 -67.39 ;
        RECT -30.73 -67.72 -30.63 -67.62 ;
        RECT -30.73 -67.95 -30.63 -67.85 ;
        RECT -30.73 -68.18 -30.63 -68.08 ;
        RECT -30.73 -68.41 -30.63 -68.31 ;
        RECT -30.73 -68.64 -30.63 -68.54 ;
        RECT 40.37 3.58 40.47 3.68 ;
        RECT 40.37 1.565 40.47 1.665 ;
        RECT 40.37 -1.665 40.47 -1.565 ;
        RECT 40.37 -4.895 40.47 -4.795 ;
        RECT 40.37 -8.125 40.47 -8.025 ;
        RECT 40.37 -11.355 40.47 -11.255 ;
        RECT 40.37 -14.585 40.47 -14.485 ;
        RECT 40.37 -17.815 40.47 -17.715 ;
        RECT 40.37 -21.045 40.47 -20.945 ;
        RECT 40.37 -24.275 40.47 -24.175 ;
        RECT 40.37 -27.505 40.47 -27.405 ;
        RECT 40.37 -30.735 40.47 -30.635 ;
        RECT 40.37 -33.965 40.47 -33.865 ;
        RECT 40.37 -37.195 40.47 -37.095 ;
        RECT 40.37 -40.425 40.47 -40.325 ;
        RECT 40.37 -43.655 40.47 -43.555 ;
        RECT 40.37 -46.885 40.47 -46.785 ;
        RECT 40.37 -50.115 40.47 -50.015 ;
        RECT 40.37 -61.015 40.47 -60.915 ;
        RECT 40.37 -66.11 40.47 -66.01 ;
        RECT 40.37 -66.34 40.47 -66.24 ;
        RECT 40.37 -66.57 40.47 -66.47 ;
        RECT 40.37 -66.8 40.47 -66.7 ;
        RECT 40.37 -67.03 40.47 -66.93 ;
        RECT 40.37 -67.26 40.47 -67.16 ;
        RECT 40.37 -67.49 40.47 -67.39 ;
        RECT 40.37 -67.72 40.47 -67.62 ;
        RECT 40.37 -67.95 40.47 -67.85 ;
        RECT 40.37 -68.18 40.47 -68.08 ;
        RECT 40.37 -68.41 40.47 -68.31 ;
        RECT 40.37 -68.64 40.47 -68.54 ;
        RECT 40.6 3.58 40.7 3.68 ;
        RECT 40.6 1.565 40.7 1.665 ;
        RECT 40.6 -1.665 40.7 -1.565 ;
        RECT 40.6 -4.895 40.7 -4.795 ;
        RECT 40.6 -8.125 40.7 -8.025 ;
        RECT 40.6 -11.355 40.7 -11.255 ;
        RECT 40.6 -14.585 40.7 -14.485 ;
        RECT 40.6 -17.815 40.7 -17.715 ;
        RECT 40.6 -21.045 40.7 -20.945 ;
        RECT 40.6 -24.275 40.7 -24.175 ;
        RECT 40.6 -27.505 40.7 -27.405 ;
        RECT 40.6 -30.735 40.7 -30.635 ;
        RECT 40.6 -33.965 40.7 -33.865 ;
        RECT 40.6 -37.195 40.7 -37.095 ;
        RECT 40.6 -40.425 40.7 -40.325 ;
        RECT 40.6 -43.655 40.7 -43.555 ;
        RECT 40.6 -46.885 40.7 -46.785 ;
        RECT 40.6 -50.115 40.7 -50.015 ;
        RECT 40.6 -61.015 40.7 -60.915 ;
        RECT 40.6 -66.11 40.7 -66.01 ;
        RECT 40.6 -66.34 40.7 -66.24 ;
        RECT 40.6 -66.57 40.7 -66.47 ;
        RECT 40.6 -66.8 40.7 -66.7 ;
        RECT 40.6 -67.03 40.7 -66.93 ;
        RECT 40.6 -67.26 40.7 -67.16 ;
        RECT 40.6 -67.49 40.7 -67.39 ;
        RECT 40.6 -67.72 40.7 -67.62 ;
        RECT 40.6 -67.95 40.7 -67.85 ;
        RECT 40.6 -68.18 40.7 -68.08 ;
        RECT 40.6 -68.41 40.7 -68.31 ;
        RECT 40.6 -68.64 40.7 -68.54 ;
        RECT 40.83 3.58 40.93 3.68 ;
        RECT 40.83 1.565 40.93 1.665 ;
        RECT 40.83 -1.665 40.93 -1.565 ;
        RECT 40.83 -4.895 40.93 -4.795 ;
        RECT 40.83 -8.125 40.93 -8.025 ;
        RECT 40.83 -11.355 40.93 -11.255 ;
        RECT 40.83 -14.585 40.93 -14.485 ;
        RECT 40.83 -17.815 40.93 -17.715 ;
        RECT 40.83 -21.045 40.93 -20.945 ;
        RECT 40.83 -24.275 40.93 -24.175 ;
        RECT 40.83 -27.505 40.93 -27.405 ;
        RECT 40.83 -30.735 40.93 -30.635 ;
        RECT 40.83 -33.965 40.93 -33.865 ;
        RECT 40.83 -37.195 40.93 -37.095 ;
        RECT 40.83 -40.425 40.93 -40.325 ;
        RECT 40.83 -43.655 40.93 -43.555 ;
        RECT 40.83 -46.885 40.93 -46.785 ;
        RECT 40.83 -50.115 40.93 -50.015 ;
        RECT 40.83 -61.015 40.93 -60.915 ;
        RECT 40.83 -66.11 40.93 -66.01 ;
        RECT 40.83 -66.34 40.93 -66.24 ;
        RECT 40.83 -66.57 40.93 -66.47 ;
        RECT 40.83 -66.8 40.93 -66.7 ;
        RECT 40.83 -67.03 40.93 -66.93 ;
        RECT 40.83 -67.26 40.93 -67.16 ;
        RECT 40.83 -67.49 40.93 -67.39 ;
        RECT 40.83 -67.72 40.93 -67.62 ;
        RECT 40.83 -67.95 40.93 -67.85 ;
        RECT 40.83 -68.18 40.93 -68.08 ;
        RECT 40.83 -68.41 40.93 -68.31 ;
        RECT 40.83 -68.64 40.93 -68.54 ;
        RECT 41.06 3.58 41.16 3.68 ;
        RECT 41.06 1.565 41.16 1.665 ;
        RECT 41.06 -1.665 41.16 -1.565 ;
        RECT 41.06 -4.895 41.16 -4.795 ;
        RECT 41.06 -8.125 41.16 -8.025 ;
        RECT 41.06 -11.355 41.16 -11.255 ;
        RECT 41.06 -14.585 41.16 -14.485 ;
        RECT 41.06 -17.815 41.16 -17.715 ;
        RECT 41.06 -21.045 41.16 -20.945 ;
        RECT 41.06 -24.275 41.16 -24.175 ;
        RECT 41.06 -27.505 41.16 -27.405 ;
        RECT 41.06 -30.735 41.16 -30.635 ;
        RECT 41.06 -33.965 41.16 -33.865 ;
        RECT 41.06 -37.195 41.16 -37.095 ;
        RECT 41.06 -40.425 41.16 -40.325 ;
        RECT 41.06 -43.655 41.16 -43.555 ;
        RECT 41.06 -46.885 41.16 -46.785 ;
        RECT 41.06 -50.115 41.16 -50.015 ;
        RECT 41.06 -61.015 41.16 -60.915 ;
        RECT 41.06 -66.11 41.16 -66.01 ;
        RECT 41.06 -66.34 41.16 -66.24 ;
        RECT 41.06 -66.57 41.16 -66.47 ;
        RECT 41.06 -66.8 41.16 -66.7 ;
        RECT 41.06 -67.03 41.16 -66.93 ;
        RECT 41.06 -67.26 41.16 -67.16 ;
        RECT 41.06 -67.49 41.16 -67.39 ;
        RECT 41.06 -67.72 41.16 -67.62 ;
        RECT 41.06 -67.95 41.16 -67.85 ;
        RECT 41.06 -68.18 41.16 -68.08 ;
        RECT 41.06 -68.41 41.16 -68.31 ;
        RECT 41.06 -68.64 41.16 -68.54 ;
    END
  END vdd!
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M1 ;
        RECT -6.655 3.435 -5.665 3.535 ;
    END
  END clk
  PIN addr4
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -29.565 -49.035 -29.385 0.645 ;
        RECT -29.565 -49.035 -29.465 3.005 ;
      LAYER M1 ;
        RECT -29.865 -47.255 -6.74 -47.155 ;
        RECT -29.865 -40.055 -6.74 -39.955 ;
        RECT -29.865 -34.335 -6.74 -34.235 ;
        RECT -29.865 -27.135 -6.74 -27.035 ;
        RECT -29.645 2.825 -29.26 3.005 ;
      LAYER V1 ;
        RECT -29.565 2.865 -29.465 2.965 ;
        RECT -29.525 -27.135 -29.425 -27.035 ;
        RECT -29.525 -34.335 -29.425 -34.235 ;
        RECT -29.525 -40.055 -29.425 -39.955 ;
        RECT -29.525 -47.255 -29.425 -47.155 ;
    END
  END addr4
  PIN addr3
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -28.965 -49.035 -28.785 0.645 ;
        RECT -28.965 -49.035 -28.865 3.345 ;
      LAYER M1 ;
        RECT -29.865 -47.475 -9.08 -47.375 ;
        RECT -29.865 -39.835 -9.08 -39.735 ;
        RECT -29.865 -21.635 -9.08 -21.535 ;
        RECT -29.865 -13.995 -9.08 -13.895 ;
        RECT -29.645 3.165 -28.66 3.345 ;
      LAYER V1 ;
        RECT -28.965 3.205 -28.865 3.305 ;
        RECT -28.925 -13.995 -28.825 -13.895 ;
        RECT -28.925 -21.635 -28.825 -21.535 ;
        RECT -28.925 -39.835 -28.825 -39.735 ;
        RECT -28.925 -47.475 -28.825 -47.375 ;
    END
  END addr3
  PIN addr2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -28.365 -49.035 -28.185 0.645 ;
        RECT -28.365 -49.035 -28.265 3.685 ;
      LAYER M1 ;
        RECT -29.865 -47.695 -9.34 -47.595 ;
        RECT -29.865 -34.775 -9.34 -34.675 ;
        RECT -29.865 -21.855 -9.34 -21.755 ;
        RECT -29.865 -8.935 -9.34 -8.835 ;
        RECT -29.645 3.505 -28.06 3.685 ;
      LAYER V1 ;
        RECT -28.365 3.545 -28.265 3.645 ;
        RECT -28.325 -8.935 -28.225 -8.835 ;
        RECT -28.325 -21.855 -28.225 -21.755 ;
        RECT -28.325 -34.775 -28.225 -34.675 ;
        RECT -28.325 -47.695 -28.225 -47.595 ;
    END
  END addr2
  PIN addr1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -27.765 -49.035 -27.585 0.645 ;
        RECT -27.765 -49.035 -27.665 4.025 ;
      LAYER M1 ;
        RECT -29.865 -47.915 -10.38 -47.815 ;
        RECT -29.865 -39.395 -10.38 -39.295 ;
        RECT -29.865 -34.995 -10.38 -34.895 ;
        RECT -29.865 -26.475 -10.38 -26.375 ;
        RECT -29.865 -22.075 -10.38 -21.975 ;
        RECT -29.865 -13.555 -10.38 -13.455 ;
        RECT -29.865 -9.155 -10.38 -9.055 ;
        RECT -29.865 -0.635 -10.38 -0.535 ;
        RECT -29.645 3.845 -27.46 4.025 ;
      LAYER V1 ;
        RECT -27.765 3.885 -27.665 3.985 ;
        RECT -27.725 -0.635 -27.625 -0.535 ;
        RECT -27.725 -9.155 -27.625 -9.055 ;
        RECT -27.725 -13.555 -27.625 -13.455 ;
        RECT -27.725 -22.075 -27.625 -21.975 ;
        RECT -27.725 -26.475 -27.625 -26.375 ;
        RECT -27.725 -34.995 -27.625 -34.895 ;
        RECT -27.725 -39.395 -27.625 -39.295 ;
        RECT -27.725 -47.915 -27.625 -47.815 ;
    END
  END addr1
  PIN addr0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -27.165 -49.035 -26.985 0.645 ;
        RECT -27.165 -49.035 -27.065 4.365 ;
      LAYER M1 ;
        RECT -29.865 -48.355 -10.64 -48.255 ;
        RECT -29.865 -38.955 -10.64 -38.855 ;
        RECT -29.865 -35.435 -10.64 -35.335 ;
        RECT -29.865 -26.035 -10.64 -25.935 ;
        RECT -29.865 -22.515 -10.64 -22.415 ;
        RECT -29.865 -13.115 -10.64 -13.015 ;
        RECT -29.865 -9.595 -10.64 -9.495 ;
        RECT -29.865 -0.195 -10.64 -0.095 ;
        RECT -29.645 4.185 -26.86 4.365 ;
      LAYER V1 ;
        RECT -27.165 4.225 -27.065 4.325 ;
        RECT -27.125 -0.195 -27.025 -0.095 ;
        RECT -27.125 -9.595 -27.025 -9.495 ;
        RECT -27.125 -13.115 -27.025 -13.015 ;
        RECT -27.125 -22.515 -27.025 -22.415 ;
        RECT -27.125 -26.035 -27.025 -25.935 ;
        RECT -27.125 -35.435 -27.025 -35.335 ;
        RECT -27.125 -38.955 -27.025 -38.855 ;
        RECT -27.125 -48.355 -27.025 -48.255 ;
    END
  END addr0
  PIN addr6
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -12.165 -55.495 -11.985 -51.035 ;
        RECT -12.165 -58.295 -12.065 -51.035 ;
      LAYER M1 ;
        RECT -12.465 -52.315 -6.48 -52.215 ;
        RECT -12.245 -58.295 -11.86 -58.115 ;
      LAYER V1 ;
        RECT -12.165 -58.255 -12.065 -58.155 ;
        RECT -12.125 -52.315 -12.025 -52.215 ;
    END
  END addr6
  PIN addr5
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -11.565 -55.495 -11.385 -51.035 ;
        RECT -11.565 -57.955 -11.465 -51.035 ;
      LAYER M1 ;
        RECT -12.465 -51.875 -6.74 -51.775 ;
        RECT -12.245 -57.955 -11.26 -57.775 ;
      LAYER V1 ;
        RECT -11.565 -57.915 -11.465 -57.815 ;
        RECT -11.525 -51.875 -11.425 -51.775 ;
    END
  END addr5
  OBS
    LAYER M1 ;
      RECT -4.705 -48.8 -4.525 -48.62 ;
      RECT -4.705 -48.755 38.5 -48.665 ;
      RECT -3.405 -48.28 -3.225 -48.1 ;
      RECT -3.405 -48.235 38.5 -48.145 ;
      RECT -2.105 -45.57 -1.925 -45.39 ;
      RECT -2.105 -45.525 38.5 -45.435 ;
      RECT -0.805 -45.05 -0.625 -44.87 ;
      RECT -0.805 -45.005 38.5 -44.915 ;
      RECT -0.805 -42.34 -0.625 -42.16 ;
      RECT -0.805 -42.295 38.5 -42.205 ;
      RECT -2.105 -41.82 -1.925 -41.64 ;
      RECT -2.105 -41.775 38.5 -41.685 ;
      RECT -3.405 -39.11 -3.225 -38.93 ;
      RECT -3.405 -39.065 38.5 -38.975 ;
      RECT -4.705 -38.59 -4.525 -38.41 ;
      RECT -4.705 -38.545 38.5 -38.455 ;
      RECT -4.705 -35.88 -4.525 -35.7 ;
      RECT -4.705 -35.835 38.5 -35.745 ;
      RECT -3.405 -35.36 -3.225 -35.18 ;
      RECT -3.405 -35.315 38.5 -35.225 ;
      RECT -2.105 -32.65 -1.925 -32.47 ;
      RECT -2.105 -32.605 38.5 -32.515 ;
      RECT -0.805 -32.13 -0.625 -31.95 ;
      RECT -0.805 -32.085 38.5 -31.995 ;
      RECT -0.805 -29.42 -0.625 -29.24 ;
      RECT -0.805 -29.375 38.5 -29.285 ;
      RECT -2.105 -28.9 -1.925 -28.72 ;
      RECT -2.105 -28.855 38.5 -28.765 ;
      RECT -3.405 -26.19 -3.225 -26.01 ;
      RECT -3.405 -26.145 38.5 -26.055 ;
      RECT -4.705 -25.67 -4.525 -25.49 ;
      RECT -4.705 -25.625 38.5 -25.535 ;
      RECT -4.705 -22.96 -4.525 -22.78 ;
      RECT -4.705 -22.915 38.5 -22.825 ;
      RECT -3.405 -22.44 -3.225 -22.26 ;
      RECT -3.405 -22.395 38.5 -22.305 ;
      RECT -2.105 -19.73 -1.925 -19.55 ;
      RECT -2.105 -19.685 38.5 -19.595 ;
      RECT -0.805 -19.21 -0.625 -19.03 ;
      RECT -0.805 -19.165 38.5 -19.075 ;
      RECT -0.805 -16.5 -0.625 -16.32 ;
      RECT -0.805 -16.455 38.5 -16.365 ;
      RECT -2.105 -15.98 -1.925 -15.8 ;
      RECT -2.105 -15.935 38.5 -15.845 ;
      RECT -3.405 -13.27 -3.225 -13.09 ;
      RECT -3.405 -13.225 38.5 -13.135 ;
      RECT -4.705 -12.75 -4.525 -12.57 ;
      RECT -4.705 -12.705 38.5 -12.615 ;
      RECT -4.705 -10.04 -4.525 -9.86 ;
      RECT -4.705 -9.995 38.5 -9.905 ;
      RECT -3.405 -9.52 -3.225 -9.34 ;
      RECT -3.405 -9.475 38.5 -9.385 ;
      RECT -2.105 -6.81 -1.925 -6.63 ;
      RECT -2.105 -6.765 38.5 -6.675 ;
      RECT -0.805 -6.29 -0.625 -6.11 ;
      RECT -0.805 -6.245 38.5 -6.155 ;
      RECT -0.805 -3.58 -0.625 -3.4 ;
      RECT -0.805 -3.535 38.5 -3.445 ;
      RECT -2.105 -3.06 -1.925 -2.88 ;
      RECT -2.105 -3.015 38.5 -2.925 ;
      RECT -3.405 -0.35 -3.225 -0.17 ;
      RECT -3.405 -0.305 38.5 -0.215 ;
      RECT -4.705 0.17 -4.525 0.35 ;
      RECT -4.705 0.215 38.5 0.305 ;
      RECT 34.635 -57.255 38.415 -57.135 ;
      RECT 35.955 -57.795 36.055 -57.135 ;
      RECT 35.395 -57.795 35.495 -57.135 ;
      RECT 34.835 -57.795 34.935 -57.135 ;
      RECT -4.705 -51.51 -4.525 -51.33 ;
      RECT -4.705 -51.465 38.28 -51.375 ;
      RECT 38.005 -49.858 38.095 -48.85 ;
      RECT 37.955 -49.255 38.095 -49.085 ;
      RECT 38.005 -48.05 38.095 -47.042 ;
      RECT 37.955 -47.815 38.095 -47.645 ;
      RECT 38.005 -46.628 38.095 -45.62 ;
      RECT 37.955 -46.025 38.095 -45.855 ;
      RECT 38.005 -44.82 38.095 -43.812 ;
      RECT 37.955 -44.585 38.095 -44.415 ;
      RECT 38.005 -43.398 38.095 -42.39 ;
      RECT 37.955 -42.795 38.095 -42.625 ;
      RECT 38.005 -41.59 38.095 -40.582 ;
      RECT 37.955 -41.355 38.095 -41.185 ;
      RECT 38.005 -40.168 38.095 -39.16 ;
      RECT 37.955 -39.565 38.095 -39.395 ;
      RECT 38.005 -38.36 38.095 -37.352 ;
      RECT 37.955 -38.125 38.095 -37.955 ;
      RECT 38.005 -36.938 38.095 -35.93 ;
      RECT 37.955 -36.335 38.095 -36.165 ;
      RECT 38.005 -35.13 38.095 -34.122 ;
      RECT 37.955 -34.895 38.095 -34.725 ;
      RECT 38.005 -33.708 38.095 -32.7 ;
      RECT 37.955 -33.105 38.095 -32.935 ;
      RECT 38.005 -31.9 38.095 -30.892 ;
      RECT 37.955 -31.665 38.095 -31.495 ;
      RECT 38.005 -30.478 38.095 -29.47 ;
      RECT 37.955 -29.875 38.095 -29.705 ;
      RECT 38.005 -28.67 38.095 -27.662 ;
      RECT 37.955 -28.435 38.095 -28.265 ;
      RECT 38.005 -27.248 38.095 -26.24 ;
      RECT 37.955 -26.645 38.095 -26.475 ;
      RECT 38.005 -25.44 38.095 -24.432 ;
      RECT 37.955 -25.205 38.095 -25.035 ;
      RECT 38.005 -24.018 38.095 -23.01 ;
      RECT 37.955 -23.415 38.095 -23.245 ;
      RECT 38.005 -22.21 38.095 -21.202 ;
      RECT 37.955 -21.975 38.095 -21.805 ;
      RECT 38.005 -20.788 38.095 -19.78 ;
      RECT 37.955 -20.185 38.095 -20.015 ;
      RECT 38.005 -18.98 38.095 -17.972 ;
      RECT 37.955 -18.745 38.095 -18.575 ;
      RECT 38.005 -17.558 38.095 -16.55 ;
      RECT 37.955 -16.955 38.095 -16.785 ;
      RECT 38.005 -15.75 38.095 -14.742 ;
      RECT 37.955 -15.515 38.095 -15.345 ;
      RECT 38.005 -14.328 38.095 -13.32 ;
      RECT 37.955 -13.725 38.095 -13.555 ;
      RECT 38.005 -12.52 38.095 -11.512 ;
      RECT 37.955 -12.285 38.095 -12.115 ;
      RECT 38.005 -11.098 38.095 -10.09 ;
      RECT 37.955 -10.495 38.095 -10.325 ;
      RECT 38.005 -9.29 38.095 -8.282 ;
      RECT 37.955 -9.055 38.095 -8.885 ;
      RECT 38.005 -7.868 38.095 -6.86 ;
      RECT 37.955 -7.265 38.095 -7.095 ;
      RECT 38.005 -6.06 38.095 -5.052 ;
      RECT 37.955 -5.825 38.095 -5.655 ;
      RECT 38.005 -4.638 38.095 -3.63 ;
      RECT 37.955 -4.035 38.095 -3.865 ;
      RECT 38.005 -2.83 38.095 -1.822 ;
      RECT 37.955 -2.595 38.095 -2.425 ;
      RECT 38.005 -1.408 38.095 -0.4 ;
      RECT 37.955 -0.805 38.095 -0.635 ;
      RECT 38.005 0.4 38.095 1.408 ;
      RECT 37.955 0.635 38.095 0.805 ;
      RECT 36.575 -60.005 38.055 -59.905 ;
      RECT 36.575 -60.515 36.675 -59.905 ;
      RECT 36.795 -57.47 38.055 -57.37 ;
      RECT 37.955 -57.795 38.055 -57.37 ;
      RECT 37.395 -57.795 37.495 -57.37 ;
      RECT 36.835 -57.795 36.935 -57.37 ;
      RECT 37.605 -49.858 37.695 -48.851 ;
      RECT 37.605 -49.545 37.745 -49.375 ;
      RECT 37.605 -48.049 37.695 -47.042 ;
      RECT 37.605 -47.525 37.745 -47.355 ;
      RECT 37.605 -46.628 37.695 -45.621 ;
      RECT 37.605 -46.315 37.745 -46.145 ;
      RECT 37.605 -44.819 37.695 -43.812 ;
      RECT 37.605 -44.295 37.745 -44.125 ;
      RECT 37.605 -43.398 37.695 -42.391 ;
      RECT 37.605 -43.085 37.745 -42.915 ;
      RECT 37.605 -41.589 37.695 -40.582 ;
      RECT 37.605 -41.065 37.745 -40.895 ;
      RECT 37.605 -40.168 37.695 -39.161 ;
      RECT 37.605 -39.855 37.745 -39.685 ;
      RECT 37.605 -38.359 37.695 -37.352 ;
      RECT 37.605 -37.835 37.745 -37.665 ;
      RECT 37.605 -36.938 37.695 -35.931 ;
      RECT 37.605 -36.625 37.745 -36.455 ;
      RECT 37.605 -35.129 37.695 -34.122 ;
      RECT 37.605 -34.605 37.745 -34.435 ;
      RECT 37.605 -33.708 37.695 -32.701 ;
      RECT 37.605 -33.395 37.745 -33.225 ;
      RECT 37.605 -31.899 37.695 -30.892 ;
      RECT 37.605 -31.375 37.745 -31.205 ;
      RECT 37.605 -30.478 37.695 -29.471 ;
      RECT 37.605 -30.165 37.745 -29.995 ;
      RECT 37.605 -28.669 37.695 -27.662 ;
      RECT 37.605 -28.145 37.745 -27.975 ;
      RECT 37.605 -27.248 37.695 -26.241 ;
      RECT 37.605 -26.935 37.745 -26.765 ;
      RECT 37.605 -25.439 37.695 -24.432 ;
      RECT 37.605 -24.915 37.745 -24.745 ;
      RECT 37.605 -24.018 37.695 -23.011 ;
      RECT 37.605 -23.705 37.745 -23.535 ;
      RECT 37.605 -22.209 37.695 -21.202 ;
      RECT 37.605 -21.685 37.745 -21.515 ;
      RECT 37.605 -20.788 37.695 -19.781 ;
      RECT 37.605 -20.475 37.745 -20.305 ;
      RECT 37.605 -18.979 37.695 -17.972 ;
      RECT 37.605 -18.455 37.745 -18.285 ;
      RECT 37.605 -17.558 37.695 -16.551 ;
      RECT 37.605 -17.245 37.745 -17.075 ;
      RECT 37.605 -15.749 37.695 -14.742 ;
      RECT 37.605 -15.225 37.745 -15.055 ;
      RECT 37.605 -14.328 37.695 -13.321 ;
      RECT 37.605 -14.015 37.745 -13.845 ;
      RECT 37.605 -12.519 37.695 -11.512 ;
      RECT 37.605 -11.995 37.745 -11.825 ;
      RECT 37.605 -11.098 37.695 -10.091 ;
      RECT 37.605 -10.785 37.745 -10.615 ;
      RECT 37.605 -9.289 37.695 -8.282 ;
      RECT 37.605 -8.765 37.745 -8.595 ;
      RECT 37.605 -7.868 37.695 -6.861 ;
      RECT 37.605 -7.555 37.745 -7.385 ;
      RECT 37.605 -6.059 37.695 -5.052 ;
      RECT 37.605 -5.535 37.745 -5.365 ;
      RECT 37.605 -4.638 37.695 -3.631 ;
      RECT 37.605 -4.325 37.745 -4.155 ;
      RECT 37.605 -2.829 37.695 -1.822 ;
      RECT 37.605 -2.305 37.745 -2.135 ;
      RECT 37.605 -1.408 37.695 -0.401 ;
      RECT 37.605 -1.095 37.745 -0.925 ;
      RECT 37.605 0.401 37.695 1.408 ;
      RECT 37.605 0.925 37.745 1.095 ;
      RECT 36.935 -59.815 37.105 -59.705 ;
      RECT 33.785 -59.815 37.105 -59.715 ;
      RECT -3.405 -52.03 -3.225 -51.85 ;
      RECT -3.405 -51.985 37.08 -51.895 ;
      RECT 36.805 -49.858 36.895 -48.85 ;
      RECT 36.755 -49.255 36.895 -49.085 ;
      RECT 36.805 -48.05 36.895 -47.042 ;
      RECT 36.755 -47.815 36.895 -47.645 ;
      RECT 36.805 -46.628 36.895 -45.62 ;
      RECT 36.755 -46.025 36.895 -45.855 ;
      RECT 36.805 -44.82 36.895 -43.812 ;
      RECT 36.755 -44.585 36.895 -44.415 ;
      RECT 36.805 -43.398 36.895 -42.39 ;
      RECT 36.755 -42.795 36.895 -42.625 ;
      RECT 36.805 -41.59 36.895 -40.582 ;
      RECT 36.755 -41.355 36.895 -41.185 ;
      RECT 36.805 -40.168 36.895 -39.16 ;
      RECT 36.755 -39.565 36.895 -39.395 ;
      RECT 36.805 -38.36 36.895 -37.352 ;
      RECT 36.755 -38.125 36.895 -37.955 ;
      RECT 36.805 -36.938 36.895 -35.93 ;
      RECT 36.755 -36.335 36.895 -36.165 ;
      RECT 36.805 -35.13 36.895 -34.122 ;
      RECT 36.755 -34.895 36.895 -34.725 ;
      RECT 36.805 -33.708 36.895 -32.7 ;
      RECT 36.755 -33.105 36.895 -32.935 ;
      RECT 36.805 -31.9 36.895 -30.892 ;
      RECT 36.755 -31.665 36.895 -31.495 ;
      RECT 36.805 -30.478 36.895 -29.47 ;
      RECT 36.755 -29.875 36.895 -29.705 ;
      RECT 36.805 -28.67 36.895 -27.662 ;
      RECT 36.755 -28.435 36.895 -28.265 ;
      RECT 36.805 -27.248 36.895 -26.24 ;
      RECT 36.755 -26.645 36.895 -26.475 ;
      RECT 36.805 -25.44 36.895 -24.432 ;
      RECT 36.755 -25.205 36.895 -25.035 ;
      RECT 36.805 -24.018 36.895 -23.01 ;
      RECT 36.755 -23.415 36.895 -23.245 ;
      RECT 36.805 -22.21 36.895 -21.202 ;
      RECT 36.755 -21.975 36.895 -21.805 ;
      RECT 36.805 -20.788 36.895 -19.78 ;
      RECT 36.755 -20.185 36.895 -20.015 ;
      RECT 36.805 -18.98 36.895 -17.972 ;
      RECT 36.755 -18.745 36.895 -18.575 ;
      RECT 36.805 -17.558 36.895 -16.55 ;
      RECT 36.755 -16.955 36.895 -16.785 ;
      RECT 36.805 -15.75 36.895 -14.742 ;
      RECT 36.755 -15.515 36.895 -15.345 ;
      RECT 36.805 -14.328 36.895 -13.32 ;
      RECT 36.755 -13.725 36.895 -13.555 ;
      RECT 36.805 -12.52 36.895 -11.512 ;
      RECT 36.755 -12.285 36.895 -12.115 ;
      RECT 36.805 -11.098 36.895 -10.09 ;
      RECT 36.755 -10.495 36.895 -10.325 ;
      RECT 36.805 -9.29 36.895 -8.282 ;
      RECT 36.755 -9.055 36.895 -8.885 ;
      RECT 36.805 -7.868 36.895 -6.86 ;
      RECT 36.755 -7.265 36.895 -7.095 ;
      RECT 36.805 -6.06 36.895 -5.052 ;
      RECT 36.755 -5.825 36.895 -5.655 ;
      RECT 36.805 -4.638 36.895 -3.63 ;
      RECT 36.755 -4.035 36.895 -3.865 ;
      RECT 36.805 -2.83 36.895 -1.822 ;
      RECT 36.755 -2.595 36.895 -2.425 ;
      RECT 36.805 -1.408 36.895 -0.4 ;
      RECT 36.755 -0.805 36.895 -0.635 ;
      RECT 36.805 0.4 36.895 1.408 ;
      RECT 36.755 0.635 36.895 0.805 ;
      RECT 36.405 -49.858 36.495 -48.851 ;
      RECT 36.405 -49.545 36.545 -49.375 ;
      RECT 36.405 -48.049 36.495 -47.042 ;
      RECT 36.405 -47.525 36.545 -47.355 ;
      RECT 36.405 -46.628 36.495 -45.621 ;
      RECT 36.405 -46.315 36.545 -46.145 ;
      RECT 36.405 -44.819 36.495 -43.812 ;
      RECT 36.405 -44.295 36.545 -44.125 ;
      RECT 36.405 -43.398 36.495 -42.391 ;
      RECT 36.405 -43.085 36.545 -42.915 ;
      RECT 36.405 -41.589 36.495 -40.582 ;
      RECT 36.405 -41.065 36.545 -40.895 ;
      RECT 36.405 -40.168 36.495 -39.161 ;
      RECT 36.405 -39.855 36.545 -39.685 ;
      RECT 36.405 -38.359 36.495 -37.352 ;
      RECT 36.405 -37.835 36.545 -37.665 ;
      RECT 36.405 -36.938 36.495 -35.931 ;
      RECT 36.405 -36.625 36.545 -36.455 ;
      RECT 36.405 -35.129 36.495 -34.122 ;
      RECT 36.405 -34.605 36.545 -34.435 ;
      RECT 36.405 -33.708 36.495 -32.701 ;
      RECT 36.405 -33.395 36.545 -33.225 ;
      RECT 36.405 -31.899 36.495 -30.892 ;
      RECT 36.405 -31.375 36.545 -31.205 ;
      RECT 36.405 -30.478 36.495 -29.471 ;
      RECT 36.405 -30.165 36.545 -29.995 ;
      RECT 36.405 -28.669 36.495 -27.662 ;
      RECT 36.405 -28.145 36.545 -27.975 ;
      RECT 36.405 -27.248 36.495 -26.241 ;
      RECT 36.405 -26.935 36.545 -26.765 ;
      RECT 36.405 -25.439 36.495 -24.432 ;
      RECT 36.405 -24.915 36.545 -24.745 ;
      RECT 36.405 -24.018 36.495 -23.011 ;
      RECT 36.405 -23.705 36.545 -23.535 ;
      RECT 36.405 -22.209 36.495 -21.202 ;
      RECT 36.405 -21.685 36.545 -21.515 ;
      RECT 36.405 -20.788 36.495 -19.781 ;
      RECT 36.405 -20.475 36.545 -20.305 ;
      RECT 36.405 -18.979 36.495 -17.972 ;
      RECT 36.405 -18.455 36.545 -18.285 ;
      RECT 36.405 -17.558 36.495 -16.551 ;
      RECT 36.405 -17.245 36.545 -17.075 ;
      RECT 36.405 -15.749 36.495 -14.742 ;
      RECT 36.405 -15.225 36.545 -15.055 ;
      RECT 36.405 -14.328 36.495 -13.321 ;
      RECT 36.405 -14.015 36.545 -13.845 ;
      RECT 36.405 -12.519 36.495 -11.512 ;
      RECT 36.405 -11.995 36.545 -11.825 ;
      RECT 36.405 -11.098 36.495 -10.091 ;
      RECT 36.405 -10.785 36.545 -10.615 ;
      RECT 36.405 -9.289 36.495 -8.282 ;
      RECT 36.405 -8.765 36.545 -8.595 ;
      RECT 36.405 -7.868 36.495 -6.861 ;
      RECT 36.405 -7.555 36.545 -7.385 ;
      RECT 36.405 -6.059 36.495 -5.052 ;
      RECT 36.405 -5.535 36.545 -5.365 ;
      RECT 36.405 -4.638 36.495 -3.631 ;
      RECT 36.405 -4.325 36.545 -4.155 ;
      RECT 36.405 -2.829 36.495 -1.822 ;
      RECT 36.405 -2.305 36.545 -2.135 ;
      RECT 36.405 -1.408 36.495 -0.401 ;
      RECT 36.405 -1.095 36.545 -0.925 ;
      RECT 36.405 0.401 36.495 1.408 ;
      RECT 36.405 0.925 36.545 1.095 ;
      RECT -4.965 -59.31 -4.785 -59.13 ;
      RECT -4.965 -59.265 36.515 -59.175 ;
      RECT 34.555 -60.005 36.035 -59.905 ;
      RECT 34.555 -60.375 34.655 -59.905 ;
      RECT 34.36 -62.715 35.935 -62.595 ;
      RECT 35.835 -63.215 35.935 -62.595 ;
      RECT 35.24 -63.215 35.34 -62.595 ;
      RECT 34.36 -63.17 34.46 -62.595 ;
      RECT -2.105 -54.74 -1.925 -54.56 ;
      RECT -2.105 -54.695 35.88 -54.605 ;
      RECT 35.605 -49.858 35.695 -48.85 ;
      RECT 35.555 -49.255 35.695 -49.085 ;
      RECT 35.605 -48.05 35.695 -47.042 ;
      RECT 35.555 -47.815 35.695 -47.645 ;
      RECT 35.605 -46.628 35.695 -45.62 ;
      RECT 35.555 -46.025 35.695 -45.855 ;
      RECT 35.605 -44.82 35.695 -43.812 ;
      RECT 35.555 -44.585 35.695 -44.415 ;
      RECT 35.605 -43.398 35.695 -42.39 ;
      RECT 35.555 -42.795 35.695 -42.625 ;
      RECT 35.605 -41.59 35.695 -40.582 ;
      RECT 35.555 -41.355 35.695 -41.185 ;
      RECT 35.605 -40.168 35.695 -39.16 ;
      RECT 35.555 -39.565 35.695 -39.395 ;
      RECT 35.605 -38.36 35.695 -37.352 ;
      RECT 35.555 -38.125 35.695 -37.955 ;
      RECT 35.605 -36.938 35.695 -35.93 ;
      RECT 35.555 -36.335 35.695 -36.165 ;
      RECT 35.605 -35.13 35.695 -34.122 ;
      RECT 35.555 -34.895 35.695 -34.725 ;
      RECT 35.605 -33.708 35.695 -32.7 ;
      RECT 35.555 -33.105 35.695 -32.935 ;
      RECT 35.605 -31.9 35.695 -30.892 ;
      RECT 35.555 -31.665 35.695 -31.495 ;
      RECT 35.605 -30.478 35.695 -29.47 ;
      RECT 35.555 -29.875 35.695 -29.705 ;
      RECT 35.605 -28.67 35.695 -27.662 ;
      RECT 35.555 -28.435 35.695 -28.265 ;
      RECT 35.605 -27.248 35.695 -26.24 ;
      RECT 35.555 -26.645 35.695 -26.475 ;
      RECT 35.605 -25.44 35.695 -24.432 ;
      RECT 35.555 -25.205 35.695 -25.035 ;
      RECT 35.605 -24.018 35.695 -23.01 ;
      RECT 35.555 -23.415 35.695 -23.245 ;
      RECT 35.605 -22.21 35.695 -21.202 ;
      RECT 35.555 -21.975 35.695 -21.805 ;
      RECT 35.605 -20.788 35.695 -19.78 ;
      RECT 35.555 -20.185 35.695 -20.015 ;
      RECT 35.605 -18.98 35.695 -17.972 ;
      RECT 35.555 -18.745 35.695 -18.575 ;
      RECT 35.605 -17.558 35.695 -16.55 ;
      RECT 35.555 -16.955 35.695 -16.785 ;
      RECT 35.605 -15.75 35.695 -14.742 ;
      RECT 35.555 -15.515 35.695 -15.345 ;
      RECT 35.605 -14.328 35.695 -13.32 ;
      RECT 35.555 -13.725 35.695 -13.555 ;
      RECT 35.605 -12.52 35.695 -11.512 ;
      RECT 35.555 -12.285 35.695 -12.115 ;
      RECT 35.605 -11.098 35.695 -10.09 ;
      RECT 35.555 -10.495 35.695 -10.325 ;
      RECT 35.605 -9.29 35.695 -8.282 ;
      RECT 35.555 -9.055 35.695 -8.885 ;
      RECT 35.605 -7.868 35.695 -6.86 ;
      RECT 35.555 -7.265 35.695 -7.095 ;
      RECT 35.605 -6.06 35.695 -5.052 ;
      RECT 35.555 -5.825 35.695 -5.655 ;
      RECT 35.605 -4.638 35.695 -3.63 ;
      RECT 35.555 -4.035 35.695 -3.865 ;
      RECT 35.605 -2.83 35.695 -1.822 ;
      RECT 35.555 -2.595 35.695 -2.425 ;
      RECT 35.605 -1.408 35.695 -0.4 ;
      RECT 35.555 -0.805 35.695 -0.635 ;
      RECT 35.605 0.4 35.695 1.408 ;
      RECT 35.555 0.635 35.695 0.805 ;
      RECT 35.48 -63.005 35.655 -62.835 ;
      RECT 35.555 -63.215 35.655 -62.835 ;
      RECT 34.595 -61.875 34.695 -61.41 ;
      RECT 34.96 -61.875 35.06 -61.42 ;
      RECT 34.595 -61.875 35.44 -61.705 ;
      RECT 35.205 -49.858 35.295 -48.851 ;
      RECT 35.205 -49.545 35.345 -49.375 ;
      RECT 35.205 -48.049 35.295 -47.042 ;
      RECT 35.205 -47.525 35.345 -47.355 ;
      RECT 35.205 -46.628 35.295 -45.621 ;
      RECT 35.205 -46.315 35.345 -46.145 ;
      RECT 35.205 -44.819 35.295 -43.812 ;
      RECT 35.205 -44.295 35.345 -44.125 ;
      RECT 35.205 -43.398 35.295 -42.391 ;
      RECT 35.205 -43.085 35.345 -42.915 ;
      RECT 35.205 -41.589 35.295 -40.582 ;
      RECT 35.205 -41.065 35.345 -40.895 ;
      RECT 35.205 -40.168 35.295 -39.161 ;
      RECT 35.205 -39.855 35.345 -39.685 ;
      RECT 35.205 -38.359 35.295 -37.352 ;
      RECT 35.205 -37.835 35.345 -37.665 ;
      RECT 35.205 -36.938 35.295 -35.931 ;
      RECT 35.205 -36.625 35.345 -36.455 ;
      RECT 35.205 -35.129 35.295 -34.122 ;
      RECT 35.205 -34.605 35.345 -34.435 ;
      RECT 35.205 -33.708 35.295 -32.701 ;
      RECT 35.205 -33.395 35.345 -33.225 ;
      RECT 35.205 -31.899 35.295 -30.892 ;
      RECT 35.205 -31.375 35.345 -31.205 ;
      RECT 35.205 -30.478 35.295 -29.471 ;
      RECT 35.205 -30.165 35.345 -29.995 ;
      RECT 35.205 -28.669 35.295 -27.662 ;
      RECT 35.205 -28.145 35.345 -27.975 ;
      RECT 35.205 -27.248 35.295 -26.241 ;
      RECT 35.205 -26.935 35.345 -26.765 ;
      RECT 35.205 -25.439 35.295 -24.432 ;
      RECT 35.205 -24.915 35.345 -24.745 ;
      RECT 35.205 -24.018 35.295 -23.011 ;
      RECT 35.205 -23.705 35.345 -23.535 ;
      RECT 35.205 -22.209 35.295 -21.202 ;
      RECT 35.205 -21.685 35.345 -21.515 ;
      RECT 35.205 -20.788 35.295 -19.781 ;
      RECT 35.205 -20.475 35.345 -20.305 ;
      RECT 35.205 -18.979 35.295 -17.972 ;
      RECT 35.205 -18.455 35.345 -18.285 ;
      RECT 35.205 -17.558 35.295 -16.551 ;
      RECT 35.205 -17.245 35.345 -17.075 ;
      RECT 35.205 -15.749 35.295 -14.742 ;
      RECT 35.205 -15.225 35.345 -15.055 ;
      RECT 35.205 -14.328 35.295 -13.321 ;
      RECT 35.205 -14.015 35.345 -13.845 ;
      RECT 35.205 -12.519 35.295 -11.512 ;
      RECT 35.205 -11.995 35.345 -11.825 ;
      RECT 35.205 -11.098 35.295 -10.091 ;
      RECT 35.205 -10.785 35.345 -10.615 ;
      RECT 35.205 -9.289 35.295 -8.282 ;
      RECT 35.205 -8.765 35.345 -8.595 ;
      RECT 35.205 -7.868 35.295 -6.861 ;
      RECT 35.205 -7.555 35.345 -7.385 ;
      RECT 35.205 -6.059 35.295 -5.052 ;
      RECT 35.205 -5.535 35.345 -5.365 ;
      RECT 35.205 -4.638 35.295 -3.631 ;
      RECT 35.205 -4.325 35.345 -4.155 ;
      RECT 35.205 -2.829 35.295 -1.822 ;
      RECT 35.205 -2.305 35.345 -2.135 ;
      RECT 35.205 -1.408 35.295 -0.401 ;
      RECT 35.205 -1.095 35.345 -0.925 ;
      RECT 35.205 0.401 35.295 1.408 ;
      RECT 35.205 0.925 35.345 1.095 ;
      RECT 34.89 -63.005 35.06 -62.835 ;
      RECT 34.96 -63.215 35.06 -62.835 ;
      RECT -0.805 -55.26 -0.625 -55.08 ;
      RECT -1.875 -55.215 34.68 -55.125 ;
      RECT 34.405 -49.858 34.495 -48.85 ;
      RECT 34.355 -49.255 34.495 -49.085 ;
      RECT 34.405 -48.05 34.495 -47.042 ;
      RECT 34.355 -47.815 34.495 -47.645 ;
      RECT 34.405 -46.628 34.495 -45.62 ;
      RECT 34.355 -46.025 34.495 -45.855 ;
      RECT 34.405 -44.82 34.495 -43.812 ;
      RECT 34.355 -44.585 34.495 -44.415 ;
      RECT 34.405 -43.398 34.495 -42.39 ;
      RECT 34.355 -42.795 34.495 -42.625 ;
      RECT 34.405 -41.59 34.495 -40.582 ;
      RECT 34.355 -41.355 34.495 -41.185 ;
      RECT 34.405 -40.168 34.495 -39.16 ;
      RECT 34.355 -39.565 34.495 -39.395 ;
      RECT 34.405 -38.36 34.495 -37.352 ;
      RECT 34.355 -38.125 34.495 -37.955 ;
      RECT 34.405 -36.938 34.495 -35.93 ;
      RECT 34.355 -36.335 34.495 -36.165 ;
      RECT 34.405 -35.13 34.495 -34.122 ;
      RECT 34.355 -34.895 34.495 -34.725 ;
      RECT 34.405 -33.708 34.495 -32.7 ;
      RECT 34.355 -33.105 34.495 -32.935 ;
      RECT 34.405 -31.9 34.495 -30.892 ;
      RECT 34.355 -31.665 34.495 -31.495 ;
      RECT 34.405 -30.478 34.495 -29.47 ;
      RECT 34.355 -29.875 34.495 -29.705 ;
      RECT 34.405 -28.67 34.495 -27.662 ;
      RECT 34.355 -28.435 34.495 -28.265 ;
      RECT 34.405 -27.248 34.495 -26.24 ;
      RECT 34.355 -26.645 34.495 -26.475 ;
      RECT 34.405 -25.44 34.495 -24.432 ;
      RECT 34.355 -25.205 34.495 -25.035 ;
      RECT 34.405 -24.018 34.495 -23.01 ;
      RECT 34.355 -23.415 34.495 -23.245 ;
      RECT 34.405 -22.21 34.495 -21.202 ;
      RECT 34.355 -21.975 34.495 -21.805 ;
      RECT 34.405 -20.788 34.495 -19.78 ;
      RECT 34.355 -20.185 34.495 -20.015 ;
      RECT 34.405 -18.98 34.495 -17.972 ;
      RECT 34.355 -18.745 34.495 -18.575 ;
      RECT 34.405 -17.558 34.495 -16.55 ;
      RECT 34.355 -16.955 34.495 -16.785 ;
      RECT 34.405 -15.75 34.495 -14.742 ;
      RECT 34.355 -15.515 34.495 -15.345 ;
      RECT 34.405 -14.328 34.495 -13.32 ;
      RECT 34.355 -13.725 34.495 -13.555 ;
      RECT 34.405 -12.52 34.495 -11.512 ;
      RECT 34.355 -12.285 34.495 -12.115 ;
      RECT 34.405 -11.098 34.495 -10.09 ;
      RECT 34.355 -10.495 34.495 -10.325 ;
      RECT 34.405 -9.29 34.495 -8.282 ;
      RECT 34.355 -9.055 34.495 -8.885 ;
      RECT 34.405 -7.868 34.495 -6.86 ;
      RECT 34.355 -7.265 34.495 -7.095 ;
      RECT 34.405 -6.06 34.495 -5.052 ;
      RECT 34.355 -5.825 34.495 -5.655 ;
      RECT 34.405 -4.638 34.495 -3.63 ;
      RECT 34.355 -4.035 34.495 -3.865 ;
      RECT 34.405 -2.83 34.495 -1.822 ;
      RECT 34.355 -2.595 34.495 -2.425 ;
      RECT 34.405 -1.408 34.495 -0.4 ;
      RECT 34.355 -0.805 34.495 -0.635 ;
      RECT 34.405 0.4 34.495 1.408 ;
      RECT 34.355 0.635 34.495 0.805 ;
      RECT 34.005 -49.858 34.095 -48.851 ;
      RECT 34.005 -49.545 34.145 -49.375 ;
      RECT 34.005 -48.049 34.095 -47.042 ;
      RECT 34.005 -47.525 34.145 -47.355 ;
      RECT 34.005 -46.628 34.095 -45.621 ;
      RECT 34.005 -46.315 34.145 -46.145 ;
      RECT 34.005 -44.819 34.095 -43.812 ;
      RECT 34.005 -44.295 34.145 -44.125 ;
      RECT 34.005 -43.398 34.095 -42.391 ;
      RECT 34.005 -43.085 34.145 -42.915 ;
      RECT 34.005 -41.589 34.095 -40.582 ;
      RECT 34.005 -41.065 34.145 -40.895 ;
      RECT 34.005 -40.168 34.095 -39.161 ;
      RECT 34.005 -39.855 34.145 -39.685 ;
      RECT 34.005 -38.359 34.095 -37.352 ;
      RECT 34.005 -37.835 34.145 -37.665 ;
      RECT 34.005 -36.938 34.095 -35.931 ;
      RECT 34.005 -36.625 34.145 -36.455 ;
      RECT 34.005 -35.129 34.095 -34.122 ;
      RECT 34.005 -34.605 34.145 -34.435 ;
      RECT 34.005 -33.708 34.095 -32.701 ;
      RECT 34.005 -33.395 34.145 -33.225 ;
      RECT 34.005 -31.899 34.095 -30.892 ;
      RECT 34.005 -31.375 34.145 -31.205 ;
      RECT 34.005 -30.478 34.095 -29.471 ;
      RECT 34.005 -30.165 34.145 -29.995 ;
      RECT 34.005 -28.669 34.095 -27.662 ;
      RECT 34.005 -28.145 34.145 -27.975 ;
      RECT 34.005 -27.248 34.095 -26.241 ;
      RECT 34.005 -26.935 34.145 -26.765 ;
      RECT 34.005 -25.439 34.095 -24.432 ;
      RECT 34.005 -24.915 34.145 -24.745 ;
      RECT 34.005 -24.018 34.095 -23.011 ;
      RECT 34.005 -23.705 34.145 -23.535 ;
      RECT 34.005 -22.209 34.095 -21.202 ;
      RECT 34.005 -21.685 34.145 -21.515 ;
      RECT 34.005 -20.788 34.095 -19.781 ;
      RECT 34.005 -20.475 34.145 -20.305 ;
      RECT 34.005 -18.979 34.095 -17.972 ;
      RECT 34.005 -18.455 34.145 -18.285 ;
      RECT 34.005 -17.558 34.095 -16.551 ;
      RECT 34.005 -17.245 34.145 -17.075 ;
      RECT 34.005 -15.749 34.095 -14.742 ;
      RECT 34.005 -15.225 34.145 -15.055 ;
      RECT 34.005 -14.328 34.095 -13.321 ;
      RECT 34.005 -14.015 34.145 -13.845 ;
      RECT 34.005 -12.519 34.095 -11.512 ;
      RECT 34.005 -11.995 34.145 -11.825 ;
      RECT 34.005 -11.098 34.095 -10.091 ;
      RECT 34.005 -10.785 34.145 -10.615 ;
      RECT 34.005 -9.289 34.095 -8.282 ;
      RECT 34.005 -8.765 34.145 -8.595 ;
      RECT 34.005 -7.868 34.095 -6.861 ;
      RECT 34.005 -7.555 34.145 -7.385 ;
      RECT 34.005 -6.059 34.095 -5.052 ;
      RECT 34.005 -5.535 34.145 -5.365 ;
      RECT 34.005 -4.638 34.095 -3.631 ;
      RECT 34.005 -4.325 34.145 -4.155 ;
      RECT 34.005 -2.829 34.095 -1.822 ;
      RECT 34.005 -2.305 34.145 -2.135 ;
      RECT 34.005 -1.408 34.095 -0.401 ;
      RECT 34.005 -1.095 34.145 -0.925 ;
      RECT 34.005 0.401 34.095 1.408 ;
      RECT 34.005 0.925 34.145 1.095 ;
      RECT 29.835 -57.255 33.615 -57.135 ;
      RECT 31.155 -57.795 31.255 -57.135 ;
      RECT 30.595 -57.795 30.695 -57.135 ;
      RECT 30.035 -57.795 30.135 -57.135 ;
      RECT 33.205 -49.858 33.295 -48.85 ;
      RECT 33.155 -49.255 33.295 -49.085 ;
      RECT 33.205 -48.05 33.295 -47.042 ;
      RECT 33.155 -47.815 33.295 -47.645 ;
      RECT 33.205 -46.628 33.295 -45.62 ;
      RECT 33.155 -46.025 33.295 -45.855 ;
      RECT 33.205 -44.82 33.295 -43.812 ;
      RECT 33.155 -44.585 33.295 -44.415 ;
      RECT 33.205 -43.398 33.295 -42.39 ;
      RECT 33.155 -42.795 33.295 -42.625 ;
      RECT 33.205 -41.59 33.295 -40.582 ;
      RECT 33.155 -41.355 33.295 -41.185 ;
      RECT 33.205 -40.168 33.295 -39.16 ;
      RECT 33.155 -39.565 33.295 -39.395 ;
      RECT 33.205 -38.36 33.295 -37.352 ;
      RECT 33.155 -38.125 33.295 -37.955 ;
      RECT 33.205 -36.938 33.295 -35.93 ;
      RECT 33.155 -36.335 33.295 -36.165 ;
      RECT 33.205 -35.13 33.295 -34.122 ;
      RECT 33.155 -34.895 33.295 -34.725 ;
      RECT 33.205 -33.708 33.295 -32.7 ;
      RECT 33.155 -33.105 33.295 -32.935 ;
      RECT 33.205 -31.9 33.295 -30.892 ;
      RECT 33.155 -31.665 33.295 -31.495 ;
      RECT 33.205 -30.478 33.295 -29.47 ;
      RECT 33.155 -29.875 33.295 -29.705 ;
      RECT 33.205 -28.67 33.295 -27.662 ;
      RECT 33.155 -28.435 33.295 -28.265 ;
      RECT 33.205 -27.248 33.295 -26.24 ;
      RECT 33.155 -26.645 33.295 -26.475 ;
      RECT 33.205 -25.44 33.295 -24.432 ;
      RECT 33.155 -25.205 33.295 -25.035 ;
      RECT 33.205 -24.018 33.295 -23.01 ;
      RECT 33.155 -23.415 33.295 -23.245 ;
      RECT 33.205 -22.21 33.295 -21.202 ;
      RECT 33.155 -21.975 33.295 -21.805 ;
      RECT 33.205 -20.788 33.295 -19.78 ;
      RECT 33.155 -20.185 33.295 -20.015 ;
      RECT 33.205 -18.98 33.295 -17.972 ;
      RECT 33.155 -18.745 33.295 -18.575 ;
      RECT 33.205 -17.558 33.295 -16.55 ;
      RECT 33.155 -16.955 33.295 -16.785 ;
      RECT 33.205 -15.75 33.295 -14.742 ;
      RECT 33.155 -15.515 33.295 -15.345 ;
      RECT 33.205 -14.328 33.295 -13.32 ;
      RECT 33.155 -13.725 33.295 -13.555 ;
      RECT 33.205 -12.52 33.295 -11.512 ;
      RECT 33.155 -12.285 33.295 -12.115 ;
      RECT 33.205 -11.098 33.295 -10.09 ;
      RECT 33.155 -10.495 33.295 -10.325 ;
      RECT 33.205 -9.29 33.295 -8.282 ;
      RECT 33.155 -9.055 33.295 -8.885 ;
      RECT 33.205 -7.868 33.295 -6.86 ;
      RECT 33.155 -7.265 33.295 -7.095 ;
      RECT 33.205 -6.06 33.295 -5.052 ;
      RECT 33.155 -5.825 33.295 -5.655 ;
      RECT 33.205 -4.638 33.295 -3.63 ;
      RECT 33.155 -4.035 33.295 -3.865 ;
      RECT 33.205 -2.83 33.295 -1.822 ;
      RECT 33.155 -2.595 33.295 -2.425 ;
      RECT 33.205 -1.408 33.295 -0.4 ;
      RECT 33.155 -0.805 33.295 -0.635 ;
      RECT 33.205 0.4 33.295 1.408 ;
      RECT 33.155 0.635 33.295 0.805 ;
      RECT 31.775 -60.005 33.255 -59.905 ;
      RECT 31.775 -60.515 31.875 -59.905 ;
      RECT 31.995 -57.47 33.255 -57.37 ;
      RECT 33.155 -57.795 33.255 -57.37 ;
      RECT 32.595 -57.795 32.695 -57.37 ;
      RECT 32.035 -57.795 32.135 -57.37 ;
      RECT 32.805 -49.858 32.895 -48.851 ;
      RECT 32.805 -49.545 32.945 -49.375 ;
      RECT 32.805 -48.049 32.895 -47.042 ;
      RECT 32.805 -47.525 32.945 -47.355 ;
      RECT 32.805 -46.628 32.895 -45.621 ;
      RECT 32.805 -46.315 32.945 -46.145 ;
      RECT 32.805 -44.819 32.895 -43.812 ;
      RECT 32.805 -44.295 32.945 -44.125 ;
      RECT 32.805 -43.398 32.895 -42.391 ;
      RECT 32.805 -43.085 32.945 -42.915 ;
      RECT 32.805 -41.589 32.895 -40.582 ;
      RECT 32.805 -41.065 32.945 -40.895 ;
      RECT 32.805 -40.168 32.895 -39.161 ;
      RECT 32.805 -39.855 32.945 -39.685 ;
      RECT 32.805 -38.359 32.895 -37.352 ;
      RECT 32.805 -37.835 32.945 -37.665 ;
      RECT 32.805 -36.938 32.895 -35.931 ;
      RECT 32.805 -36.625 32.945 -36.455 ;
      RECT 32.805 -35.129 32.895 -34.122 ;
      RECT 32.805 -34.605 32.945 -34.435 ;
      RECT 32.805 -33.708 32.895 -32.701 ;
      RECT 32.805 -33.395 32.945 -33.225 ;
      RECT 32.805 -31.899 32.895 -30.892 ;
      RECT 32.805 -31.375 32.945 -31.205 ;
      RECT 32.805 -30.478 32.895 -29.471 ;
      RECT 32.805 -30.165 32.945 -29.995 ;
      RECT 32.805 -28.669 32.895 -27.662 ;
      RECT 32.805 -28.145 32.945 -27.975 ;
      RECT 32.805 -27.248 32.895 -26.241 ;
      RECT 32.805 -26.935 32.945 -26.765 ;
      RECT 32.805 -25.439 32.895 -24.432 ;
      RECT 32.805 -24.915 32.945 -24.745 ;
      RECT 32.805 -24.018 32.895 -23.011 ;
      RECT 32.805 -23.705 32.945 -23.535 ;
      RECT 32.805 -22.209 32.895 -21.202 ;
      RECT 32.805 -21.685 32.945 -21.515 ;
      RECT 32.805 -20.788 32.895 -19.781 ;
      RECT 32.805 -20.475 32.945 -20.305 ;
      RECT 32.805 -18.979 32.895 -17.972 ;
      RECT 32.805 -18.455 32.945 -18.285 ;
      RECT 32.805 -17.558 32.895 -16.551 ;
      RECT 32.805 -17.245 32.945 -17.075 ;
      RECT 32.805 -15.749 32.895 -14.742 ;
      RECT 32.805 -15.225 32.945 -15.055 ;
      RECT 32.805 -14.328 32.895 -13.321 ;
      RECT 32.805 -14.015 32.945 -13.845 ;
      RECT 32.805 -12.519 32.895 -11.512 ;
      RECT 32.805 -11.995 32.945 -11.825 ;
      RECT 32.805 -11.098 32.895 -10.091 ;
      RECT 32.805 -10.785 32.945 -10.615 ;
      RECT 32.805 -9.289 32.895 -8.282 ;
      RECT 32.805 -8.765 32.945 -8.595 ;
      RECT 32.805 -7.868 32.895 -6.861 ;
      RECT 32.805 -7.555 32.945 -7.385 ;
      RECT 32.805 -6.059 32.895 -5.052 ;
      RECT 32.805 -5.535 32.945 -5.365 ;
      RECT 32.805 -4.638 32.895 -3.631 ;
      RECT 32.805 -4.325 32.945 -4.155 ;
      RECT 32.805 -2.829 32.895 -1.822 ;
      RECT 32.805 -2.305 32.945 -2.135 ;
      RECT 32.805 -1.408 32.895 -0.401 ;
      RECT 32.805 -1.095 32.945 -0.925 ;
      RECT 32.805 0.401 32.895 1.408 ;
      RECT 32.805 0.925 32.945 1.095 ;
      RECT 32.135 -59.815 32.305 -59.705 ;
      RECT 28.985 -59.815 32.305 -59.715 ;
      RECT 32.005 -49.858 32.095 -48.85 ;
      RECT 31.955 -49.255 32.095 -49.085 ;
      RECT 32.005 -48.05 32.095 -47.042 ;
      RECT 31.955 -47.815 32.095 -47.645 ;
      RECT 32.005 -46.628 32.095 -45.62 ;
      RECT 31.955 -46.025 32.095 -45.855 ;
      RECT 32.005 -44.82 32.095 -43.812 ;
      RECT 31.955 -44.585 32.095 -44.415 ;
      RECT 32.005 -43.398 32.095 -42.39 ;
      RECT 31.955 -42.795 32.095 -42.625 ;
      RECT 32.005 -41.59 32.095 -40.582 ;
      RECT 31.955 -41.355 32.095 -41.185 ;
      RECT 32.005 -40.168 32.095 -39.16 ;
      RECT 31.955 -39.565 32.095 -39.395 ;
      RECT 32.005 -38.36 32.095 -37.352 ;
      RECT 31.955 -38.125 32.095 -37.955 ;
      RECT 32.005 -36.938 32.095 -35.93 ;
      RECT 31.955 -36.335 32.095 -36.165 ;
      RECT 32.005 -35.13 32.095 -34.122 ;
      RECT 31.955 -34.895 32.095 -34.725 ;
      RECT 32.005 -33.708 32.095 -32.7 ;
      RECT 31.955 -33.105 32.095 -32.935 ;
      RECT 32.005 -31.9 32.095 -30.892 ;
      RECT 31.955 -31.665 32.095 -31.495 ;
      RECT 32.005 -30.478 32.095 -29.47 ;
      RECT 31.955 -29.875 32.095 -29.705 ;
      RECT 32.005 -28.67 32.095 -27.662 ;
      RECT 31.955 -28.435 32.095 -28.265 ;
      RECT 32.005 -27.248 32.095 -26.24 ;
      RECT 31.955 -26.645 32.095 -26.475 ;
      RECT 32.005 -25.44 32.095 -24.432 ;
      RECT 31.955 -25.205 32.095 -25.035 ;
      RECT 32.005 -24.018 32.095 -23.01 ;
      RECT 31.955 -23.415 32.095 -23.245 ;
      RECT 32.005 -22.21 32.095 -21.202 ;
      RECT 31.955 -21.975 32.095 -21.805 ;
      RECT 32.005 -20.788 32.095 -19.78 ;
      RECT 31.955 -20.185 32.095 -20.015 ;
      RECT 32.005 -18.98 32.095 -17.972 ;
      RECT 31.955 -18.745 32.095 -18.575 ;
      RECT 32.005 -17.558 32.095 -16.55 ;
      RECT 31.955 -16.955 32.095 -16.785 ;
      RECT 32.005 -15.75 32.095 -14.742 ;
      RECT 31.955 -15.515 32.095 -15.345 ;
      RECT 32.005 -14.328 32.095 -13.32 ;
      RECT 31.955 -13.725 32.095 -13.555 ;
      RECT 32.005 -12.52 32.095 -11.512 ;
      RECT 31.955 -12.285 32.095 -12.115 ;
      RECT 32.005 -11.098 32.095 -10.09 ;
      RECT 31.955 -10.495 32.095 -10.325 ;
      RECT 32.005 -9.29 32.095 -8.282 ;
      RECT 31.955 -9.055 32.095 -8.885 ;
      RECT 32.005 -7.868 32.095 -6.86 ;
      RECT 31.955 -7.265 32.095 -7.095 ;
      RECT 32.005 -6.06 32.095 -5.052 ;
      RECT 31.955 -5.825 32.095 -5.655 ;
      RECT 32.005 -4.638 32.095 -3.63 ;
      RECT 31.955 -4.035 32.095 -3.865 ;
      RECT 32.005 -2.83 32.095 -1.822 ;
      RECT 31.955 -2.595 32.095 -2.425 ;
      RECT 32.005 -1.408 32.095 -0.4 ;
      RECT 31.955 -0.805 32.095 -0.635 ;
      RECT 32.005 0.4 32.095 1.408 ;
      RECT 31.955 0.635 32.095 0.805 ;
      RECT 31.605 -49.858 31.695 -48.851 ;
      RECT 31.605 -49.545 31.745 -49.375 ;
      RECT 31.605 -48.049 31.695 -47.042 ;
      RECT 31.605 -47.525 31.745 -47.355 ;
      RECT 31.605 -46.628 31.695 -45.621 ;
      RECT 31.605 -46.315 31.745 -46.145 ;
      RECT 31.605 -44.819 31.695 -43.812 ;
      RECT 31.605 -44.295 31.745 -44.125 ;
      RECT 31.605 -43.398 31.695 -42.391 ;
      RECT 31.605 -43.085 31.745 -42.915 ;
      RECT 31.605 -41.589 31.695 -40.582 ;
      RECT 31.605 -41.065 31.745 -40.895 ;
      RECT 31.605 -40.168 31.695 -39.161 ;
      RECT 31.605 -39.855 31.745 -39.685 ;
      RECT 31.605 -38.359 31.695 -37.352 ;
      RECT 31.605 -37.835 31.745 -37.665 ;
      RECT 31.605 -36.938 31.695 -35.931 ;
      RECT 31.605 -36.625 31.745 -36.455 ;
      RECT 31.605 -35.129 31.695 -34.122 ;
      RECT 31.605 -34.605 31.745 -34.435 ;
      RECT 31.605 -33.708 31.695 -32.701 ;
      RECT 31.605 -33.395 31.745 -33.225 ;
      RECT 31.605 -31.899 31.695 -30.892 ;
      RECT 31.605 -31.375 31.745 -31.205 ;
      RECT 31.605 -30.478 31.695 -29.471 ;
      RECT 31.605 -30.165 31.745 -29.995 ;
      RECT 31.605 -28.669 31.695 -27.662 ;
      RECT 31.605 -28.145 31.745 -27.975 ;
      RECT 31.605 -27.248 31.695 -26.241 ;
      RECT 31.605 -26.935 31.745 -26.765 ;
      RECT 31.605 -25.439 31.695 -24.432 ;
      RECT 31.605 -24.915 31.745 -24.745 ;
      RECT 31.605 -24.018 31.695 -23.011 ;
      RECT 31.605 -23.705 31.745 -23.535 ;
      RECT 31.605 -22.209 31.695 -21.202 ;
      RECT 31.605 -21.685 31.745 -21.515 ;
      RECT 31.605 -20.788 31.695 -19.781 ;
      RECT 31.605 -20.475 31.745 -20.305 ;
      RECT 31.605 -18.979 31.695 -17.972 ;
      RECT 31.605 -18.455 31.745 -18.285 ;
      RECT 31.605 -17.558 31.695 -16.551 ;
      RECT 31.605 -17.245 31.745 -17.075 ;
      RECT 31.605 -15.749 31.695 -14.742 ;
      RECT 31.605 -15.225 31.745 -15.055 ;
      RECT 31.605 -14.328 31.695 -13.321 ;
      RECT 31.605 -14.015 31.745 -13.845 ;
      RECT 31.605 -12.519 31.695 -11.512 ;
      RECT 31.605 -11.995 31.745 -11.825 ;
      RECT 31.605 -11.098 31.695 -10.091 ;
      RECT 31.605 -10.785 31.745 -10.615 ;
      RECT 31.605 -9.289 31.695 -8.282 ;
      RECT 31.605 -8.765 31.745 -8.595 ;
      RECT 31.605 -7.868 31.695 -6.861 ;
      RECT 31.605 -7.555 31.745 -7.385 ;
      RECT 31.605 -6.059 31.695 -5.052 ;
      RECT 31.605 -5.535 31.745 -5.365 ;
      RECT 31.605 -4.638 31.695 -3.631 ;
      RECT 31.605 -4.325 31.745 -4.155 ;
      RECT 31.605 -2.829 31.695 -1.822 ;
      RECT 31.605 -2.305 31.745 -2.135 ;
      RECT 31.605 -1.408 31.695 -0.401 ;
      RECT 31.605 -1.095 31.745 -0.925 ;
      RECT 31.605 0.401 31.695 1.408 ;
      RECT 31.605 0.925 31.745 1.095 ;
      RECT 29.755 -60.005 31.235 -59.905 ;
      RECT 29.755 -60.375 29.855 -59.905 ;
      RECT 29.56 -62.715 31.135 -62.595 ;
      RECT 31.035 -63.215 31.135 -62.595 ;
      RECT 30.44 -63.215 30.54 -62.595 ;
      RECT 29.56 -63.17 29.66 -62.595 ;
      RECT 30.805 -49.858 30.895 -48.85 ;
      RECT 30.755 -49.255 30.895 -49.085 ;
      RECT 30.805 -48.05 30.895 -47.042 ;
      RECT 30.755 -47.815 30.895 -47.645 ;
      RECT 30.805 -46.628 30.895 -45.62 ;
      RECT 30.755 -46.025 30.895 -45.855 ;
      RECT 30.805 -44.82 30.895 -43.812 ;
      RECT 30.755 -44.585 30.895 -44.415 ;
      RECT 30.805 -43.398 30.895 -42.39 ;
      RECT 30.755 -42.795 30.895 -42.625 ;
      RECT 30.805 -41.59 30.895 -40.582 ;
      RECT 30.755 -41.355 30.895 -41.185 ;
      RECT 30.805 -40.168 30.895 -39.16 ;
      RECT 30.755 -39.565 30.895 -39.395 ;
      RECT 30.805 -38.36 30.895 -37.352 ;
      RECT 30.755 -38.125 30.895 -37.955 ;
      RECT 30.805 -36.938 30.895 -35.93 ;
      RECT 30.755 -36.335 30.895 -36.165 ;
      RECT 30.805 -35.13 30.895 -34.122 ;
      RECT 30.755 -34.895 30.895 -34.725 ;
      RECT 30.805 -33.708 30.895 -32.7 ;
      RECT 30.755 -33.105 30.895 -32.935 ;
      RECT 30.805 -31.9 30.895 -30.892 ;
      RECT 30.755 -31.665 30.895 -31.495 ;
      RECT 30.805 -30.478 30.895 -29.47 ;
      RECT 30.755 -29.875 30.895 -29.705 ;
      RECT 30.805 -28.67 30.895 -27.662 ;
      RECT 30.755 -28.435 30.895 -28.265 ;
      RECT 30.805 -27.248 30.895 -26.24 ;
      RECT 30.755 -26.645 30.895 -26.475 ;
      RECT 30.805 -25.44 30.895 -24.432 ;
      RECT 30.755 -25.205 30.895 -25.035 ;
      RECT 30.805 -24.018 30.895 -23.01 ;
      RECT 30.755 -23.415 30.895 -23.245 ;
      RECT 30.805 -22.21 30.895 -21.202 ;
      RECT 30.755 -21.975 30.895 -21.805 ;
      RECT 30.805 -20.788 30.895 -19.78 ;
      RECT 30.755 -20.185 30.895 -20.015 ;
      RECT 30.805 -18.98 30.895 -17.972 ;
      RECT 30.755 -18.745 30.895 -18.575 ;
      RECT 30.805 -17.558 30.895 -16.55 ;
      RECT 30.755 -16.955 30.895 -16.785 ;
      RECT 30.805 -15.75 30.895 -14.742 ;
      RECT 30.755 -15.515 30.895 -15.345 ;
      RECT 30.805 -14.328 30.895 -13.32 ;
      RECT 30.755 -13.725 30.895 -13.555 ;
      RECT 30.805 -12.52 30.895 -11.512 ;
      RECT 30.755 -12.285 30.895 -12.115 ;
      RECT 30.805 -11.098 30.895 -10.09 ;
      RECT 30.755 -10.495 30.895 -10.325 ;
      RECT 30.805 -9.29 30.895 -8.282 ;
      RECT 30.755 -9.055 30.895 -8.885 ;
      RECT 30.805 -7.868 30.895 -6.86 ;
      RECT 30.755 -7.265 30.895 -7.095 ;
      RECT 30.805 -6.06 30.895 -5.052 ;
      RECT 30.755 -5.825 30.895 -5.655 ;
      RECT 30.805 -4.638 30.895 -3.63 ;
      RECT 30.755 -4.035 30.895 -3.865 ;
      RECT 30.805 -2.83 30.895 -1.822 ;
      RECT 30.755 -2.595 30.895 -2.425 ;
      RECT 30.805 -1.408 30.895 -0.4 ;
      RECT 30.755 -0.805 30.895 -0.635 ;
      RECT 30.805 0.4 30.895 1.408 ;
      RECT 30.755 0.635 30.895 0.805 ;
      RECT 30.68 -63.005 30.855 -62.835 ;
      RECT 30.755 -63.215 30.855 -62.835 ;
      RECT 29.795 -61.875 29.895 -61.41 ;
      RECT 30.16 -61.875 30.26 -61.42 ;
      RECT 29.795 -61.875 30.64 -61.705 ;
      RECT 30.405 -49.858 30.495 -48.851 ;
      RECT 30.405 -49.545 30.545 -49.375 ;
      RECT 30.405 -48.049 30.495 -47.042 ;
      RECT 30.405 -47.525 30.545 -47.355 ;
      RECT 30.405 -46.628 30.495 -45.621 ;
      RECT 30.405 -46.315 30.545 -46.145 ;
      RECT 30.405 -44.819 30.495 -43.812 ;
      RECT 30.405 -44.295 30.545 -44.125 ;
      RECT 30.405 -43.398 30.495 -42.391 ;
      RECT 30.405 -43.085 30.545 -42.915 ;
      RECT 30.405 -41.589 30.495 -40.582 ;
      RECT 30.405 -41.065 30.545 -40.895 ;
      RECT 30.405 -40.168 30.495 -39.161 ;
      RECT 30.405 -39.855 30.545 -39.685 ;
      RECT 30.405 -38.359 30.495 -37.352 ;
      RECT 30.405 -37.835 30.545 -37.665 ;
      RECT 30.405 -36.938 30.495 -35.931 ;
      RECT 30.405 -36.625 30.545 -36.455 ;
      RECT 30.405 -35.129 30.495 -34.122 ;
      RECT 30.405 -34.605 30.545 -34.435 ;
      RECT 30.405 -33.708 30.495 -32.701 ;
      RECT 30.405 -33.395 30.545 -33.225 ;
      RECT 30.405 -31.899 30.495 -30.892 ;
      RECT 30.405 -31.375 30.545 -31.205 ;
      RECT 30.405 -30.478 30.495 -29.471 ;
      RECT 30.405 -30.165 30.545 -29.995 ;
      RECT 30.405 -28.669 30.495 -27.662 ;
      RECT 30.405 -28.145 30.545 -27.975 ;
      RECT 30.405 -27.248 30.495 -26.241 ;
      RECT 30.405 -26.935 30.545 -26.765 ;
      RECT 30.405 -25.439 30.495 -24.432 ;
      RECT 30.405 -24.915 30.545 -24.745 ;
      RECT 30.405 -24.018 30.495 -23.011 ;
      RECT 30.405 -23.705 30.545 -23.535 ;
      RECT 30.405 -22.209 30.495 -21.202 ;
      RECT 30.405 -21.685 30.545 -21.515 ;
      RECT 30.405 -20.788 30.495 -19.781 ;
      RECT 30.405 -20.475 30.545 -20.305 ;
      RECT 30.405 -18.979 30.495 -17.972 ;
      RECT 30.405 -18.455 30.545 -18.285 ;
      RECT 30.405 -17.558 30.495 -16.551 ;
      RECT 30.405 -17.245 30.545 -17.075 ;
      RECT 30.405 -15.749 30.495 -14.742 ;
      RECT 30.405 -15.225 30.545 -15.055 ;
      RECT 30.405 -14.328 30.495 -13.321 ;
      RECT 30.405 -14.015 30.545 -13.845 ;
      RECT 30.405 -12.519 30.495 -11.512 ;
      RECT 30.405 -11.995 30.545 -11.825 ;
      RECT 30.405 -11.098 30.495 -10.091 ;
      RECT 30.405 -10.785 30.545 -10.615 ;
      RECT 30.405 -9.289 30.495 -8.282 ;
      RECT 30.405 -8.765 30.545 -8.595 ;
      RECT 30.405 -7.868 30.495 -6.861 ;
      RECT 30.405 -7.555 30.545 -7.385 ;
      RECT 30.405 -6.059 30.495 -5.052 ;
      RECT 30.405 -5.535 30.545 -5.365 ;
      RECT 30.405 -4.638 30.495 -3.631 ;
      RECT 30.405 -4.325 30.545 -4.155 ;
      RECT 30.405 -2.829 30.495 -1.822 ;
      RECT 30.405 -2.305 30.545 -2.135 ;
      RECT 30.405 -1.408 30.495 -0.401 ;
      RECT 30.405 -1.095 30.545 -0.925 ;
      RECT 30.405 0.401 30.495 1.408 ;
      RECT 30.405 0.925 30.545 1.095 ;
      RECT 30.09 -63.005 30.26 -62.835 ;
      RECT 30.16 -63.215 30.26 -62.835 ;
      RECT 29.605 -49.858 29.695 -48.85 ;
      RECT 29.555 -49.255 29.695 -49.085 ;
      RECT 29.605 -48.05 29.695 -47.042 ;
      RECT 29.555 -47.815 29.695 -47.645 ;
      RECT 29.605 -46.628 29.695 -45.62 ;
      RECT 29.555 -46.025 29.695 -45.855 ;
      RECT 29.605 -44.82 29.695 -43.812 ;
      RECT 29.555 -44.585 29.695 -44.415 ;
      RECT 29.605 -43.398 29.695 -42.39 ;
      RECT 29.555 -42.795 29.695 -42.625 ;
      RECT 29.605 -41.59 29.695 -40.582 ;
      RECT 29.555 -41.355 29.695 -41.185 ;
      RECT 29.605 -40.168 29.695 -39.16 ;
      RECT 29.555 -39.565 29.695 -39.395 ;
      RECT 29.605 -38.36 29.695 -37.352 ;
      RECT 29.555 -38.125 29.695 -37.955 ;
      RECT 29.605 -36.938 29.695 -35.93 ;
      RECT 29.555 -36.335 29.695 -36.165 ;
      RECT 29.605 -35.13 29.695 -34.122 ;
      RECT 29.555 -34.895 29.695 -34.725 ;
      RECT 29.605 -33.708 29.695 -32.7 ;
      RECT 29.555 -33.105 29.695 -32.935 ;
      RECT 29.605 -31.9 29.695 -30.892 ;
      RECT 29.555 -31.665 29.695 -31.495 ;
      RECT 29.605 -30.478 29.695 -29.47 ;
      RECT 29.555 -29.875 29.695 -29.705 ;
      RECT 29.605 -28.67 29.695 -27.662 ;
      RECT 29.555 -28.435 29.695 -28.265 ;
      RECT 29.605 -27.248 29.695 -26.24 ;
      RECT 29.555 -26.645 29.695 -26.475 ;
      RECT 29.605 -25.44 29.695 -24.432 ;
      RECT 29.555 -25.205 29.695 -25.035 ;
      RECT 29.605 -24.018 29.695 -23.01 ;
      RECT 29.555 -23.415 29.695 -23.245 ;
      RECT 29.605 -22.21 29.695 -21.202 ;
      RECT 29.555 -21.975 29.695 -21.805 ;
      RECT 29.605 -20.788 29.695 -19.78 ;
      RECT 29.555 -20.185 29.695 -20.015 ;
      RECT 29.605 -18.98 29.695 -17.972 ;
      RECT 29.555 -18.745 29.695 -18.575 ;
      RECT 29.605 -17.558 29.695 -16.55 ;
      RECT 29.555 -16.955 29.695 -16.785 ;
      RECT 29.605 -15.75 29.695 -14.742 ;
      RECT 29.555 -15.515 29.695 -15.345 ;
      RECT 29.605 -14.328 29.695 -13.32 ;
      RECT 29.555 -13.725 29.695 -13.555 ;
      RECT 29.605 -12.52 29.695 -11.512 ;
      RECT 29.555 -12.285 29.695 -12.115 ;
      RECT 29.605 -11.098 29.695 -10.09 ;
      RECT 29.555 -10.495 29.695 -10.325 ;
      RECT 29.605 -9.29 29.695 -8.282 ;
      RECT 29.555 -9.055 29.695 -8.885 ;
      RECT 29.605 -7.868 29.695 -6.86 ;
      RECT 29.555 -7.265 29.695 -7.095 ;
      RECT 29.605 -6.06 29.695 -5.052 ;
      RECT 29.555 -5.825 29.695 -5.655 ;
      RECT 29.605 -4.638 29.695 -3.63 ;
      RECT 29.555 -4.035 29.695 -3.865 ;
      RECT 29.605 -2.83 29.695 -1.822 ;
      RECT 29.555 -2.595 29.695 -2.425 ;
      RECT 29.605 -1.408 29.695 -0.4 ;
      RECT 29.555 -0.805 29.695 -0.635 ;
      RECT 29.605 0.4 29.695 1.408 ;
      RECT 29.555 0.635 29.695 0.805 ;
      RECT 29.205 -49.858 29.295 -48.851 ;
      RECT 29.205 -49.545 29.345 -49.375 ;
      RECT 29.205 -48.049 29.295 -47.042 ;
      RECT 29.205 -47.525 29.345 -47.355 ;
      RECT 29.205 -46.628 29.295 -45.621 ;
      RECT 29.205 -46.315 29.345 -46.145 ;
      RECT 29.205 -44.819 29.295 -43.812 ;
      RECT 29.205 -44.295 29.345 -44.125 ;
      RECT 29.205 -43.398 29.295 -42.391 ;
      RECT 29.205 -43.085 29.345 -42.915 ;
      RECT 29.205 -41.589 29.295 -40.582 ;
      RECT 29.205 -41.065 29.345 -40.895 ;
      RECT 29.205 -40.168 29.295 -39.161 ;
      RECT 29.205 -39.855 29.345 -39.685 ;
      RECT 29.205 -38.359 29.295 -37.352 ;
      RECT 29.205 -37.835 29.345 -37.665 ;
      RECT 29.205 -36.938 29.295 -35.931 ;
      RECT 29.205 -36.625 29.345 -36.455 ;
      RECT 29.205 -35.129 29.295 -34.122 ;
      RECT 29.205 -34.605 29.345 -34.435 ;
      RECT 29.205 -33.708 29.295 -32.701 ;
      RECT 29.205 -33.395 29.345 -33.225 ;
      RECT 29.205 -31.899 29.295 -30.892 ;
      RECT 29.205 -31.375 29.345 -31.205 ;
      RECT 29.205 -30.478 29.295 -29.471 ;
      RECT 29.205 -30.165 29.345 -29.995 ;
      RECT 29.205 -28.669 29.295 -27.662 ;
      RECT 29.205 -28.145 29.345 -27.975 ;
      RECT 29.205 -27.248 29.295 -26.241 ;
      RECT 29.205 -26.935 29.345 -26.765 ;
      RECT 29.205 -25.439 29.295 -24.432 ;
      RECT 29.205 -24.915 29.345 -24.745 ;
      RECT 29.205 -24.018 29.295 -23.011 ;
      RECT 29.205 -23.705 29.345 -23.535 ;
      RECT 29.205 -22.209 29.295 -21.202 ;
      RECT 29.205 -21.685 29.345 -21.515 ;
      RECT 29.205 -20.788 29.295 -19.781 ;
      RECT 29.205 -20.475 29.345 -20.305 ;
      RECT 29.205 -18.979 29.295 -17.972 ;
      RECT 29.205 -18.455 29.345 -18.285 ;
      RECT 29.205 -17.558 29.295 -16.551 ;
      RECT 29.205 -17.245 29.345 -17.075 ;
      RECT 29.205 -15.749 29.295 -14.742 ;
      RECT 29.205 -15.225 29.345 -15.055 ;
      RECT 29.205 -14.328 29.295 -13.321 ;
      RECT 29.205 -14.015 29.345 -13.845 ;
      RECT 29.205 -12.519 29.295 -11.512 ;
      RECT 29.205 -11.995 29.345 -11.825 ;
      RECT 29.205 -11.098 29.295 -10.091 ;
      RECT 29.205 -10.785 29.345 -10.615 ;
      RECT 29.205 -9.289 29.295 -8.282 ;
      RECT 29.205 -8.765 29.345 -8.595 ;
      RECT 29.205 -7.868 29.295 -6.861 ;
      RECT 29.205 -7.555 29.345 -7.385 ;
      RECT 29.205 -6.059 29.295 -5.052 ;
      RECT 29.205 -5.535 29.345 -5.365 ;
      RECT 29.205 -4.638 29.295 -3.631 ;
      RECT 29.205 -4.325 29.345 -4.155 ;
      RECT 29.205 -2.829 29.295 -1.822 ;
      RECT 29.205 -2.305 29.345 -2.135 ;
      RECT 29.205 -1.408 29.295 -0.401 ;
      RECT 29.205 -1.095 29.345 -0.925 ;
      RECT 29.205 0.401 29.295 1.408 ;
      RECT 29.205 0.925 29.345 1.095 ;
      RECT 25.035 -57.255 28.815 -57.135 ;
      RECT 26.355 -57.795 26.455 -57.135 ;
      RECT 25.795 -57.795 25.895 -57.135 ;
      RECT 25.235 -57.795 25.335 -57.135 ;
      RECT 28.405 -49.858 28.495 -48.85 ;
      RECT 28.355 -49.255 28.495 -49.085 ;
      RECT 28.405 -48.05 28.495 -47.042 ;
      RECT 28.355 -47.815 28.495 -47.645 ;
      RECT 28.405 -46.628 28.495 -45.62 ;
      RECT 28.355 -46.025 28.495 -45.855 ;
      RECT 28.405 -44.82 28.495 -43.812 ;
      RECT 28.355 -44.585 28.495 -44.415 ;
      RECT 28.405 -43.398 28.495 -42.39 ;
      RECT 28.355 -42.795 28.495 -42.625 ;
      RECT 28.405 -41.59 28.495 -40.582 ;
      RECT 28.355 -41.355 28.495 -41.185 ;
      RECT 28.405 -40.168 28.495 -39.16 ;
      RECT 28.355 -39.565 28.495 -39.395 ;
      RECT 28.405 -38.36 28.495 -37.352 ;
      RECT 28.355 -38.125 28.495 -37.955 ;
      RECT 28.405 -36.938 28.495 -35.93 ;
      RECT 28.355 -36.335 28.495 -36.165 ;
      RECT 28.405 -35.13 28.495 -34.122 ;
      RECT 28.355 -34.895 28.495 -34.725 ;
      RECT 28.405 -33.708 28.495 -32.7 ;
      RECT 28.355 -33.105 28.495 -32.935 ;
      RECT 28.405 -31.9 28.495 -30.892 ;
      RECT 28.355 -31.665 28.495 -31.495 ;
      RECT 28.405 -30.478 28.495 -29.47 ;
      RECT 28.355 -29.875 28.495 -29.705 ;
      RECT 28.405 -28.67 28.495 -27.662 ;
      RECT 28.355 -28.435 28.495 -28.265 ;
      RECT 28.405 -27.248 28.495 -26.24 ;
      RECT 28.355 -26.645 28.495 -26.475 ;
      RECT 28.405 -25.44 28.495 -24.432 ;
      RECT 28.355 -25.205 28.495 -25.035 ;
      RECT 28.405 -24.018 28.495 -23.01 ;
      RECT 28.355 -23.415 28.495 -23.245 ;
      RECT 28.405 -22.21 28.495 -21.202 ;
      RECT 28.355 -21.975 28.495 -21.805 ;
      RECT 28.405 -20.788 28.495 -19.78 ;
      RECT 28.355 -20.185 28.495 -20.015 ;
      RECT 28.405 -18.98 28.495 -17.972 ;
      RECT 28.355 -18.745 28.495 -18.575 ;
      RECT 28.405 -17.558 28.495 -16.55 ;
      RECT 28.355 -16.955 28.495 -16.785 ;
      RECT 28.405 -15.75 28.495 -14.742 ;
      RECT 28.355 -15.515 28.495 -15.345 ;
      RECT 28.405 -14.328 28.495 -13.32 ;
      RECT 28.355 -13.725 28.495 -13.555 ;
      RECT 28.405 -12.52 28.495 -11.512 ;
      RECT 28.355 -12.285 28.495 -12.115 ;
      RECT 28.405 -11.098 28.495 -10.09 ;
      RECT 28.355 -10.495 28.495 -10.325 ;
      RECT 28.405 -9.29 28.495 -8.282 ;
      RECT 28.355 -9.055 28.495 -8.885 ;
      RECT 28.405 -7.868 28.495 -6.86 ;
      RECT 28.355 -7.265 28.495 -7.095 ;
      RECT 28.405 -6.06 28.495 -5.052 ;
      RECT 28.355 -5.825 28.495 -5.655 ;
      RECT 28.405 -4.638 28.495 -3.63 ;
      RECT 28.355 -4.035 28.495 -3.865 ;
      RECT 28.405 -2.83 28.495 -1.822 ;
      RECT 28.355 -2.595 28.495 -2.425 ;
      RECT 28.405 -1.408 28.495 -0.4 ;
      RECT 28.355 -0.805 28.495 -0.635 ;
      RECT 28.405 0.4 28.495 1.408 ;
      RECT 28.355 0.635 28.495 0.805 ;
      RECT 26.975 -60.005 28.455 -59.905 ;
      RECT 26.975 -60.515 27.075 -59.905 ;
      RECT 27.195 -57.47 28.455 -57.37 ;
      RECT 28.355 -57.795 28.455 -57.37 ;
      RECT 27.795 -57.795 27.895 -57.37 ;
      RECT 27.235 -57.795 27.335 -57.37 ;
      RECT 28.005 -49.858 28.095 -48.851 ;
      RECT 28.005 -49.545 28.145 -49.375 ;
      RECT 28.005 -48.049 28.095 -47.042 ;
      RECT 28.005 -47.525 28.145 -47.355 ;
      RECT 28.005 -46.628 28.095 -45.621 ;
      RECT 28.005 -46.315 28.145 -46.145 ;
      RECT 28.005 -44.819 28.095 -43.812 ;
      RECT 28.005 -44.295 28.145 -44.125 ;
      RECT 28.005 -43.398 28.095 -42.391 ;
      RECT 28.005 -43.085 28.145 -42.915 ;
      RECT 28.005 -41.589 28.095 -40.582 ;
      RECT 28.005 -41.065 28.145 -40.895 ;
      RECT 28.005 -40.168 28.095 -39.161 ;
      RECT 28.005 -39.855 28.145 -39.685 ;
      RECT 28.005 -38.359 28.095 -37.352 ;
      RECT 28.005 -37.835 28.145 -37.665 ;
      RECT 28.005 -36.938 28.095 -35.931 ;
      RECT 28.005 -36.625 28.145 -36.455 ;
      RECT 28.005 -35.129 28.095 -34.122 ;
      RECT 28.005 -34.605 28.145 -34.435 ;
      RECT 28.005 -33.708 28.095 -32.701 ;
      RECT 28.005 -33.395 28.145 -33.225 ;
      RECT 28.005 -31.899 28.095 -30.892 ;
      RECT 28.005 -31.375 28.145 -31.205 ;
      RECT 28.005 -30.478 28.095 -29.471 ;
      RECT 28.005 -30.165 28.145 -29.995 ;
      RECT 28.005 -28.669 28.095 -27.662 ;
      RECT 28.005 -28.145 28.145 -27.975 ;
      RECT 28.005 -27.248 28.095 -26.241 ;
      RECT 28.005 -26.935 28.145 -26.765 ;
      RECT 28.005 -25.439 28.095 -24.432 ;
      RECT 28.005 -24.915 28.145 -24.745 ;
      RECT 28.005 -24.018 28.095 -23.011 ;
      RECT 28.005 -23.705 28.145 -23.535 ;
      RECT 28.005 -22.209 28.095 -21.202 ;
      RECT 28.005 -21.685 28.145 -21.515 ;
      RECT 28.005 -20.788 28.095 -19.781 ;
      RECT 28.005 -20.475 28.145 -20.305 ;
      RECT 28.005 -18.979 28.095 -17.972 ;
      RECT 28.005 -18.455 28.145 -18.285 ;
      RECT 28.005 -17.558 28.095 -16.551 ;
      RECT 28.005 -17.245 28.145 -17.075 ;
      RECT 28.005 -15.749 28.095 -14.742 ;
      RECT 28.005 -15.225 28.145 -15.055 ;
      RECT 28.005 -14.328 28.095 -13.321 ;
      RECT 28.005 -14.015 28.145 -13.845 ;
      RECT 28.005 -12.519 28.095 -11.512 ;
      RECT 28.005 -11.995 28.145 -11.825 ;
      RECT 28.005 -11.098 28.095 -10.091 ;
      RECT 28.005 -10.785 28.145 -10.615 ;
      RECT 28.005 -9.289 28.095 -8.282 ;
      RECT 28.005 -8.765 28.145 -8.595 ;
      RECT 28.005 -7.868 28.095 -6.861 ;
      RECT 28.005 -7.555 28.145 -7.385 ;
      RECT 28.005 -6.059 28.095 -5.052 ;
      RECT 28.005 -5.535 28.145 -5.365 ;
      RECT 28.005 -4.638 28.095 -3.631 ;
      RECT 28.005 -4.325 28.145 -4.155 ;
      RECT 28.005 -2.829 28.095 -1.822 ;
      RECT 28.005 -2.305 28.145 -2.135 ;
      RECT 28.005 -1.408 28.095 -0.401 ;
      RECT 28.005 -1.095 28.145 -0.925 ;
      RECT 28.005 0.401 28.095 1.408 ;
      RECT 28.005 0.925 28.145 1.095 ;
      RECT 27.335 -59.815 27.505 -59.705 ;
      RECT 24.185 -59.815 27.505 -59.715 ;
      RECT 27.205 -49.858 27.295 -48.85 ;
      RECT 27.155 -49.255 27.295 -49.085 ;
      RECT 27.205 -48.05 27.295 -47.042 ;
      RECT 27.155 -47.815 27.295 -47.645 ;
      RECT 27.205 -46.628 27.295 -45.62 ;
      RECT 27.155 -46.025 27.295 -45.855 ;
      RECT 27.205 -44.82 27.295 -43.812 ;
      RECT 27.155 -44.585 27.295 -44.415 ;
      RECT 27.205 -43.398 27.295 -42.39 ;
      RECT 27.155 -42.795 27.295 -42.625 ;
      RECT 27.205 -41.59 27.295 -40.582 ;
      RECT 27.155 -41.355 27.295 -41.185 ;
      RECT 27.205 -40.168 27.295 -39.16 ;
      RECT 27.155 -39.565 27.295 -39.395 ;
      RECT 27.205 -38.36 27.295 -37.352 ;
      RECT 27.155 -38.125 27.295 -37.955 ;
      RECT 27.205 -36.938 27.295 -35.93 ;
      RECT 27.155 -36.335 27.295 -36.165 ;
      RECT 27.205 -35.13 27.295 -34.122 ;
      RECT 27.155 -34.895 27.295 -34.725 ;
      RECT 27.205 -33.708 27.295 -32.7 ;
      RECT 27.155 -33.105 27.295 -32.935 ;
      RECT 27.205 -31.9 27.295 -30.892 ;
      RECT 27.155 -31.665 27.295 -31.495 ;
      RECT 27.205 -30.478 27.295 -29.47 ;
      RECT 27.155 -29.875 27.295 -29.705 ;
      RECT 27.205 -28.67 27.295 -27.662 ;
      RECT 27.155 -28.435 27.295 -28.265 ;
      RECT 27.205 -27.248 27.295 -26.24 ;
      RECT 27.155 -26.645 27.295 -26.475 ;
      RECT 27.205 -25.44 27.295 -24.432 ;
      RECT 27.155 -25.205 27.295 -25.035 ;
      RECT 27.205 -24.018 27.295 -23.01 ;
      RECT 27.155 -23.415 27.295 -23.245 ;
      RECT 27.205 -22.21 27.295 -21.202 ;
      RECT 27.155 -21.975 27.295 -21.805 ;
      RECT 27.205 -20.788 27.295 -19.78 ;
      RECT 27.155 -20.185 27.295 -20.015 ;
      RECT 27.205 -18.98 27.295 -17.972 ;
      RECT 27.155 -18.745 27.295 -18.575 ;
      RECT 27.205 -17.558 27.295 -16.55 ;
      RECT 27.155 -16.955 27.295 -16.785 ;
      RECT 27.205 -15.75 27.295 -14.742 ;
      RECT 27.155 -15.515 27.295 -15.345 ;
      RECT 27.205 -14.328 27.295 -13.32 ;
      RECT 27.155 -13.725 27.295 -13.555 ;
      RECT 27.205 -12.52 27.295 -11.512 ;
      RECT 27.155 -12.285 27.295 -12.115 ;
      RECT 27.205 -11.098 27.295 -10.09 ;
      RECT 27.155 -10.495 27.295 -10.325 ;
      RECT 27.205 -9.29 27.295 -8.282 ;
      RECT 27.155 -9.055 27.295 -8.885 ;
      RECT 27.205 -7.868 27.295 -6.86 ;
      RECT 27.155 -7.265 27.295 -7.095 ;
      RECT 27.205 -6.06 27.295 -5.052 ;
      RECT 27.155 -5.825 27.295 -5.655 ;
      RECT 27.205 -4.638 27.295 -3.63 ;
      RECT 27.155 -4.035 27.295 -3.865 ;
      RECT 27.205 -2.83 27.295 -1.822 ;
      RECT 27.155 -2.595 27.295 -2.425 ;
      RECT 27.205 -1.408 27.295 -0.4 ;
      RECT 27.155 -0.805 27.295 -0.635 ;
      RECT 27.205 0.4 27.295 1.408 ;
      RECT 27.155 0.635 27.295 0.805 ;
      RECT 26.805 -49.858 26.895 -48.851 ;
      RECT 26.805 -49.545 26.945 -49.375 ;
      RECT 26.805 -48.049 26.895 -47.042 ;
      RECT 26.805 -47.525 26.945 -47.355 ;
      RECT 26.805 -46.628 26.895 -45.621 ;
      RECT 26.805 -46.315 26.945 -46.145 ;
      RECT 26.805 -44.819 26.895 -43.812 ;
      RECT 26.805 -44.295 26.945 -44.125 ;
      RECT 26.805 -43.398 26.895 -42.391 ;
      RECT 26.805 -43.085 26.945 -42.915 ;
      RECT 26.805 -41.589 26.895 -40.582 ;
      RECT 26.805 -41.065 26.945 -40.895 ;
      RECT 26.805 -40.168 26.895 -39.161 ;
      RECT 26.805 -39.855 26.945 -39.685 ;
      RECT 26.805 -38.359 26.895 -37.352 ;
      RECT 26.805 -37.835 26.945 -37.665 ;
      RECT 26.805 -36.938 26.895 -35.931 ;
      RECT 26.805 -36.625 26.945 -36.455 ;
      RECT 26.805 -35.129 26.895 -34.122 ;
      RECT 26.805 -34.605 26.945 -34.435 ;
      RECT 26.805 -33.708 26.895 -32.701 ;
      RECT 26.805 -33.395 26.945 -33.225 ;
      RECT 26.805 -31.899 26.895 -30.892 ;
      RECT 26.805 -31.375 26.945 -31.205 ;
      RECT 26.805 -30.478 26.895 -29.471 ;
      RECT 26.805 -30.165 26.945 -29.995 ;
      RECT 26.805 -28.669 26.895 -27.662 ;
      RECT 26.805 -28.145 26.945 -27.975 ;
      RECT 26.805 -27.248 26.895 -26.241 ;
      RECT 26.805 -26.935 26.945 -26.765 ;
      RECT 26.805 -25.439 26.895 -24.432 ;
      RECT 26.805 -24.915 26.945 -24.745 ;
      RECT 26.805 -24.018 26.895 -23.011 ;
      RECT 26.805 -23.705 26.945 -23.535 ;
      RECT 26.805 -22.209 26.895 -21.202 ;
      RECT 26.805 -21.685 26.945 -21.515 ;
      RECT 26.805 -20.788 26.895 -19.781 ;
      RECT 26.805 -20.475 26.945 -20.305 ;
      RECT 26.805 -18.979 26.895 -17.972 ;
      RECT 26.805 -18.455 26.945 -18.285 ;
      RECT 26.805 -17.558 26.895 -16.551 ;
      RECT 26.805 -17.245 26.945 -17.075 ;
      RECT 26.805 -15.749 26.895 -14.742 ;
      RECT 26.805 -15.225 26.945 -15.055 ;
      RECT 26.805 -14.328 26.895 -13.321 ;
      RECT 26.805 -14.015 26.945 -13.845 ;
      RECT 26.805 -12.519 26.895 -11.512 ;
      RECT 26.805 -11.995 26.945 -11.825 ;
      RECT 26.805 -11.098 26.895 -10.091 ;
      RECT 26.805 -10.785 26.945 -10.615 ;
      RECT 26.805 -9.289 26.895 -8.282 ;
      RECT 26.805 -8.765 26.945 -8.595 ;
      RECT 26.805 -7.868 26.895 -6.861 ;
      RECT 26.805 -7.555 26.945 -7.385 ;
      RECT 26.805 -6.059 26.895 -5.052 ;
      RECT 26.805 -5.535 26.945 -5.365 ;
      RECT 26.805 -4.638 26.895 -3.631 ;
      RECT 26.805 -4.325 26.945 -4.155 ;
      RECT 26.805 -2.829 26.895 -1.822 ;
      RECT 26.805 -2.305 26.945 -2.135 ;
      RECT 26.805 -1.408 26.895 -0.401 ;
      RECT 26.805 -1.095 26.945 -0.925 ;
      RECT 26.805 0.401 26.895 1.408 ;
      RECT 26.805 0.925 26.945 1.095 ;
      RECT 24.955 -60.005 26.435 -59.905 ;
      RECT 24.955 -60.375 25.055 -59.905 ;
      RECT 24.76 -62.715 26.335 -62.595 ;
      RECT 26.235 -63.215 26.335 -62.595 ;
      RECT 25.64 -63.215 25.74 -62.595 ;
      RECT 24.76 -63.17 24.86 -62.595 ;
      RECT 26.005 -49.858 26.095 -48.85 ;
      RECT 25.955 -49.255 26.095 -49.085 ;
      RECT 26.005 -48.05 26.095 -47.042 ;
      RECT 25.955 -47.815 26.095 -47.645 ;
      RECT 26.005 -46.628 26.095 -45.62 ;
      RECT 25.955 -46.025 26.095 -45.855 ;
      RECT 26.005 -44.82 26.095 -43.812 ;
      RECT 25.955 -44.585 26.095 -44.415 ;
      RECT 26.005 -43.398 26.095 -42.39 ;
      RECT 25.955 -42.795 26.095 -42.625 ;
      RECT 26.005 -41.59 26.095 -40.582 ;
      RECT 25.955 -41.355 26.095 -41.185 ;
      RECT 26.005 -40.168 26.095 -39.16 ;
      RECT 25.955 -39.565 26.095 -39.395 ;
      RECT 26.005 -38.36 26.095 -37.352 ;
      RECT 25.955 -38.125 26.095 -37.955 ;
      RECT 26.005 -36.938 26.095 -35.93 ;
      RECT 25.955 -36.335 26.095 -36.165 ;
      RECT 26.005 -35.13 26.095 -34.122 ;
      RECT 25.955 -34.895 26.095 -34.725 ;
      RECT 26.005 -33.708 26.095 -32.7 ;
      RECT 25.955 -33.105 26.095 -32.935 ;
      RECT 26.005 -31.9 26.095 -30.892 ;
      RECT 25.955 -31.665 26.095 -31.495 ;
      RECT 26.005 -30.478 26.095 -29.47 ;
      RECT 25.955 -29.875 26.095 -29.705 ;
      RECT 26.005 -28.67 26.095 -27.662 ;
      RECT 25.955 -28.435 26.095 -28.265 ;
      RECT 26.005 -27.248 26.095 -26.24 ;
      RECT 25.955 -26.645 26.095 -26.475 ;
      RECT 26.005 -25.44 26.095 -24.432 ;
      RECT 25.955 -25.205 26.095 -25.035 ;
      RECT 26.005 -24.018 26.095 -23.01 ;
      RECT 25.955 -23.415 26.095 -23.245 ;
      RECT 26.005 -22.21 26.095 -21.202 ;
      RECT 25.955 -21.975 26.095 -21.805 ;
      RECT 26.005 -20.788 26.095 -19.78 ;
      RECT 25.955 -20.185 26.095 -20.015 ;
      RECT 26.005 -18.98 26.095 -17.972 ;
      RECT 25.955 -18.745 26.095 -18.575 ;
      RECT 26.005 -17.558 26.095 -16.55 ;
      RECT 25.955 -16.955 26.095 -16.785 ;
      RECT 26.005 -15.75 26.095 -14.742 ;
      RECT 25.955 -15.515 26.095 -15.345 ;
      RECT 26.005 -14.328 26.095 -13.32 ;
      RECT 25.955 -13.725 26.095 -13.555 ;
      RECT 26.005 -12.52 26.095 -11.512 ;
      RECT 25.955 -12.285 26.095 -12.115 ;
      RECT 26.005 -11.098 26.095 -10.09 ;
      RECT 25.955 -10.495 26.095 -10.325 ;
      RECT 26.005 -9.29 26.095 -8.282 ;
      RECT 25.955 -9.055 26.095 -8.885 ;
      RECT 26.005 -7.868 26.095 -6.86 ;
      RECT 25.955 -7.265 26.095 -7.095 ;
      RECT 26.005 -6.06 26.095 -5.052 ;
      RECT 25.955 -5.825 26.095 -5.655 ;
      RECT 26.005 -4.638 26.095 -3.63 ;
      RECT 25.955 -4.035 26.095 -3.865 ;
      RECT 26.005 -2.83 26.095 -1.822 ;
      RECT 25.955 -2.595 26.095 -2.425 ;
      RECT 26.005 -1.408 26.095 -0.4 ;
      RECT 25.955 -0.805 26.095 -0.635 ;
      RECT 26.005 0.4 26.095 1.408 ;
      RECT 25.955 0.635 26.095 0.805 ;
      RECT 25.88 -63.005 26.055 -62.835 ;
      RECT 25.955 -63.215 26.055 -62.835 ;
      RECT 24.995 -61.875 25.095 -61.41 ;
      RECT 25.36 -61.875 25.46 -61.42 ;
      RECT 24.995 -61.875 25.84 -61.705 ;
      RECT 25.605 -49.858 25.695 -48.851 ;
      RECT 25.605 -49.545 25.745 -49.375 ;
      RECT 25.605 -48.049 25.695 -47.042 ;
      RECT 25.605 -47.525 25.745 -47.355 ;
      RECT 25.605 -46.628 25.695 -45.621 ;
      RECT 25.605 -46.315 25.745 -46.145 ;
      RECT 25.605 -44.819 25.695 -43.812 ;
      RECT 25.605 -44.295 25.745 -44.125 ;
      RECT 25.605 -43.398 25.695 -42.391 ;
      RECT 25.605 -43.085 25.745 -42.915 ;
      RECT 25.605 -41.589 25.695 -40.582 ;
      RECT 25.605 -41.065 25.745 -40.895 ;
      RECT 25.605 -40.168 25.695 -39.161 ;
      RECT 25.605 -39.855 25.745 -39.685 ;
      RECT 25.605 -38.359 25.695 -37.352 ;
      RECT 25.605 -37.835 25.745 -37.665 ;
      RECT 25.605 -36.938 25.695 -35.931 ;
      RECT 25.605 -36.625 25.745 -36.455 ;
      RECT 25.605 -35.129 25.695 -34.122 ;
      RECT 25.605 -34.605 25.745 -34.435 ;
      RECT 25.605 -33.708 25.695 -32.701 ;
      RECT 25.605 -33.395 25.745 -33.225 ;
      RECT 25.605 -31.899 25.695 -30.892 ;
      RECT 25.605 -31.375 25.745 -31.205 ;
      RECT 25.605 -30.478 25.695 -29.471 ;
      RECT 25.605 -30.165 25.745 -29.995 ;
      RECT 25.605 -28.669 25.695 -27.662 ;
      RECT 25.605 -28.145 25.745 -27.975 ;
      RECT 25.605 -27.248 25.695 -26.241 ;
      RECT 25.605 -26.935 25.745 -26.765 ;
      RECT 25.605 -25.439 25.695 -24.432 ;
      RECT 25.605 -24.915 25.745 -24.745 ;
      RECT 25.605 -24.018 25.695 -23.011 ;
      RECT 25.605 -23.705 25.745 -23.535 ;
      RECT 25.605 -22.209 25.695 -21.202 ;
      RECT 25.605 -21.685 25.745 -21.515 ;
      RECT 25.605 -20.788 25.695 -19.781 ;
      RECT 25.605 -20.475 25.745 -20.305 ;
      RECT 25.605 -18.979 25.695 -17.972 ;
      RECT 25.605 -18.455 25.745 -18.285 ;
      RECT 25.605 -17.558 25.695 -16.551 ;
      RECT 25.605 -17.245 25.745 -17.075 ;
      RECT 25.605 -15.749 25.695 -14.742 ;
      RECT 25.605 -15.225 25.745 -15.055 ;
      RECT 25.605 -14.328 25.695 -13.321 ;
      RECT 25.605 -14.015 25.745 -13.845 ;
      RECT 25.605 -12.519 25.695 -11.512 ;
      RECT 25.605 -11.995 25.745 -11.825 ;
      RECT 25.605 -11.098 25.695 -10.091 ;
      RECT 25.605 -10.785 25.745 -10.615 ;
      RECT 25.605 -9.289 25.695 -8.282 ;
      RECT 25.605 -8.765 25.745 -8.595 ;
      RECT 25.605 -7.868 25.695 -6.861 ;
      RECT 25.605 -7.555 25.745 -7.385 ;
      RECT 25.605 -6.059 25.695 -5.052 ;
      RECT 25.605 -5.535 25.745 -5.365 ;
      RECT 25.605 -4.638 25.695 -3.631 ;
      RECT 25.605 -4.325 25.745 -4.155 ;
      RECT 25.605 -2.829 25.695 -1.822 ;
      RECT 25.605 -2.305 25.745 -2.135 ;
      RECT 25.605 -1.408 25.695 -0.401 ;
      RECT 25.605 -1.095 25.745 -0.925 ;
      RECT 25.605 0.401 25.695 1.408 ;
      RECT 25.605 0.925 25.745 1.095 ;
      RECT 25.29 -63.005 25.46 -62.835 ;
      RECT 25.36 -63.215 25.46 -62.835 ;
      RECT 24.805 -49.858 24.895 -48.85 ;
      RECT 24.755 -49.255 24.895 -49.085 ;
      RECT 24.805 -48.05 24.895 -47.042 ;
      RECT 24.755 -47.815 24.895 -47.645 ;
      RECT 24.805 -46.628 24.895 -45.62 ;
      RECT 24.755 -46.025 24.895 -45.855 ;
      RECT 24.805 -44.82 24.895 -43.812 ;
      RECT 24.755 -44.585 24.895 -44.415 ;
      RECT 24.805 -43.398 24.895 -42.39 ;
      RECT 24.755 -42.795 24.895 -42.625 ;
      RECT 24.805 -41.59 24.895 -40.582 ;
      RECT 24.755 -41.355 24.895 -41.185 ;
      RECT 24.805 -40.168 24.895 -39.16 ;
      RECT 24.755 -39.565 24.895 -39.395 ;
      RECT 24.805 -38.36 24.895 -37.352 ;
      RECT 24.755 -38.125 24.895 -37.955 ;
      RECT 24.805 -36.938 24.895 -35.93 ;
      RECT 24.755 -36.335 24.895 -36.165 ;
      RECT 24.805 -35.13 24.895 -34.122 ;
      RECT 24.755 -34.895 24.895 -34.725 ;
      RECT 24.805 -33.708 24.895 -32.7 ;
      RECT 24.755 -33.105 24.895 -32.935 ;
      RECT 24.805 -31.9 24.895 -30.892 ;
      RECT 24.755 -31.665 24.895 -31.495 ;
      RECT 24.805 -30.478 24.895 -29.47 ;
      RECT 24.755 -29.875 24.895 -29.705 ;
      RECT 24.805 -28.67 24.895 -27.662 ;
      RECT 24.755 -28.435 24.895 -28.265 ;
      RECT 24.805 -27.248 24.895 -26.24 ;
      RECT 24.755 -26.645 24.895 -26.475 ;
      RECT 24.805 -25.44 24.895 -24.432 ;
      RECT 24.755 -25.205 24.895 -25.035 ;
      RECT 24.805 -24.018 24.895 -23.01 ;
      RECT 24.755 -23.415 24.895 -23.245 ;
      RECT 24.805 -22.21 24.895 -21.202 ;
      RECT 24.755 -21.975 24.895 -21.805 ;
      RECT 24.805 -20.788 24.895 -19.78 ;
      RECT 24.755 -20.185 24.895 -20.015 ;
      RECT 24.805 -18.98 24.895 -17.972 ;
      RECT 24.755 -18.745 24.895 -18.575 ;
      RECT 24.805 -17.558 24.895 -16.55 ;
      RECT 24.755 -16.955 24.895 -16.785 ;
      RECT 24.805 -15.75 24.895 -14.742 ;
      RECT 24.755 -15.515 24.895 -15.345 ;
      RECT 24.805 -14.328 24.895 -13.32 ;
      RECT 24.755 -13.725 24.895 -13.555 ;
      RECT 24.805 -12.52 24.895 -11.512 ;
      RECT 24.755 -12.285 24.895 -12.115 ;
      RECT 24.805 -11.098 24.895 -10.09 ;
      RECT 24.755 -10.495 24.895 -10.325 ;
      RECT 24.805 -9.29 24.895 -8.282 ;
      RECT 24.755 -9.055 24.895 -8.885 ;
      RECT 24.805 -7.868 24.895 -6.86 ;
      RECT 24.755 -7.265 24.895 -7.095 ;
      RECT 24.805 -6.06 24.895 -5.052 ;
      RECT 24.755 -5.825 24.895 -5.655 ;
      RECT 24.805 -4.638 24.895 -3.63 ;
      RECT 24.755 -4.035 24.895 -3.865 ;
      RECT 24.805 -2.83 24.895 -1.822 ;
      RECT 24.755 -2.595 24.895 -2.425 ;
      RECT 24.805 -1.408 24.895 -0.4 ;
      RECT 24.755 -0.805 24.895 -0.635 ;
      RECT 24.805 0.4 24.895 1.408 ;
      RECT 24.755 0.635 24.895 0.805 ;
      RECT 24.405 -49.858 24.495 -48.851 ;
      RECT 24.405 -49.545 24.545 -49.375 ;
      RECT 24.405 -48.049 24.495 -47.042 ;
      RECT 24.405 -47.525 24.545 -47.355 ;
      RECT 24.405 -46.628 24.495 -45.621 ;
      RECT 24.405 -46.315 24.545 -46.145 ;
      RECT 24.405 -44.819 24.495 -43.812 ;
      RECT 24.405 -44.295 24.545 -44.125 ;
      RECT 24.405 -43.398 24.495 -42.391 ;
      RECT 24.405 -43.085 24.545 -42.915 ;
      RECT 24.405 -41.589 24.495 -40.582 ;
      RECT 24.405 -41.065 24.545 -40.895 ;
      RECT 24.405 -40.168 24.495 -39.161 ;
      RECT 24.405 -39.855 24.545 -39.685 ;
      RECT 24.405 -38.359 24.495 -37.352 ;
      RECT 24.405 -37.835 24.545 -37.665 ;
      RECT 24.405 -36.938 24.495 -35.931 ;
      RECT 24.405 -36.625 24.545 -36.455 ;
      RECT 24.405 -35.129 24.495 -34.122 ;
      RECT 24.405 -34.605 24.545 -34.435 ;
      RECT 24.405 -33.708 24.495 -32.701 ;
      RECT 24.405 -33.395 24.545 -33.225 ;
      RECT 24.405 -31.899 24.495 -30.892 ;
      RECT 24.405 -31.375 24.545 -31.205 ;
      RECT 24.405 -30.478 24.495 -29.471 ;
      RECT 24.405 -30.165 24.545 -29.995 ;
      RECT 24.405 -28.669 24.495 -27.662 ;
      RECT 24.405 -28.145 24.545 -27.975 ;
      RECT 24.405 -27.248 24.495 -26.241 ;
      RECT 24.405 -26.935 24.545 -26.765 ;
      RECT 24.405 -25.439 24.495 -24.432 ;
      RECT 24.405 -24.915 24.545 -24.745 ;
      RECT 24.405 -24.018 24.495 -23.011 ;
      RECT 24.405 -23.705 24.545 -23.535 ;
      RECT 24.405 -22.209 24.495 -21.202 ;
      RECT 24.405 -21.685 24.545 -21.515 ;
      RECT 24.405 -20.788 24.495 -19.781 ;
      RECT 24.405 -20.475 24.545 -20.305 ;
      RECT 24.405 -18.979 24.495 -17.972 ;
      RECT 24.405 -18.455 24.545 -18.285 ;
      RECT 24.405 -17.558 24.495 -16.551 ;
      RECT 24.405 -17.245 24.545 -17.075 ;
      RECT 24.405 -15.749 24.495 -14.742 ;
      RECT 24.405 -15.225 24.545 -15.055 ;
      RECT 24.405 -14.328 24.495 -13.321 ;
      RECT 24.405 -14.015 24.545 -13.845 ;
      RECT 24.405 -12.519 24.495 -11.512 ;
      RECT 24.405 -11.995 24.545 -11.825 ;
      RECT 24.405 -11.098 24.495 -10.091 ;
      RECT 24.405 -10.785 24.545 -10.615 ;
      RECT 24.405 -9.289 24.495 -8.282 ;
      RECT 24.405 -8.765 24.545 -8.595 ;
      RECT 24.405 -7.868 24.495 -6.861 ;
      RECT 24.405 -7.555 24.545 -7.385 ;
      RECT 24.405 -6.059 24.495 -5.052 ;
      RECT 24.405 -5.535 24.545 -5.365 ;
      RECT 24.405 -4.638 24.495 -3.631 ;
      RECT 24.405 -4.325 24.545 -4.155 ;
      RECT 24.405 -2.829 24.495 -1.822 ;
      RECT 24.405 -2.305 24.545 -2.135 ;
      RECT 24.405 -1.408 24.495 -0.401 ;
      RECT 24.405 -1.095 24.545 -0.925 ;
      RECT 24.405 0.401 24.495 1.408 ;
      RECT 24.405 0.925 24.545 1.095 ;
      RECT 20.235 -57.255 24.015 -57.135 ;
      RECT 21.555 -57.795 21.655 -57.135 ;
      RECT 20.995 -57.795 21.095 -57.135 ;
      RECT 20.435 -57.795 20.535 -57.135 ;
      RECT 23.605 -49.858 23.695 -48.85 ;
      RECT 23.555 -49.255 23.695 -49.085 ;
      RECT 23.605 -48.05 23.695 -47.042 ;
      RECT 23.555 -47.815 23.695 -47.645 ;
      RECT 23.605 -46.628 23.695 -45.62 ;
      RECT 23.555 -46.025 23.695 -45.855 ;
      RECT 23.605 -44.82 23.695 -43.812 ;
      RECT 23.555 -44.585 23.695 -44.415 ;
      RECT 23.605 -43.398 23.695 -42.39 ;
      RECT 23.555 -42.795 23.695 -42.625 ;
      RECT 23.605 -41.59 23.695 -40.582 ;
      RECT 23.555 -41.355 23.695 -41.185 ;
      RECT 23.605 -40.168 23.695 -39.16 ;
      RECT 23.555 -39.565 23.695 -39.395 ;
      RECT 23.605 -38.36 23.695 -37.352 ;
      RECT 23.555 -38.125 23.695 -37.955 ;
      RECT 23.605 -36.938 23.695 -35.93 ;
      RECT 23.555 -36.335 23.695 -36.165 ;
      RECT 23.605 -35.13 23.695 -34.122 ;
      RECT 23.555 -34.895 23.695 -34.725 ;
      RECT 23.605 -33.708 23.695 -32.7 ;
      RECT 23.555 -33.105 23.695 -32.935 ;
      RECT 23.605 -31.9 23.695 -30.892 ;
      RECT 23.555 -31.665 23.695 -31.495 ;
      RECT 23.605 -30.478 23.695 -29.47 ;
      RECT 23.555 -29.875 23.695 -29.705 ;
      RECT 23.605 -28.67 23.695 -27.662 ;
      RECT 23.555 -28.435 23.695 -28.265 ;
      RECT 23.605 -27.248 23.695 -26.24 ;
      RECT 23.555 -26.645 23.695 -26.475 ;
      RECT 23.605 -25.44 23.695 -24.432 ;
      RECT 23.555 -25.205 23.695 -25.035 ;
      RECT 23.605 -24.018 23.695 -23.01 ;
      RECT 23.555 -23.415 23.695 -23.245 ;
      RECT 23.605 -22.21 23.695 -21.202 ;
      RECT 23.555 -21.975 23.695 -21.805 ;
      RECT 23.605 -20.788 23.695 -19.78 ;
      RECT 23.555 -20.185 23.695 -20.015 ;
      RECT 23.605 -18.98 23.695 -17.972 ;
      RECT 23.555 -18.745 23.695 -18.575 ;
      RECT 23.605 -17.558 23.695 -16.55 ;
      RECT 23.555 -16.955 23.695 -16.785 ;
      RECT 23.605 -15.75 23.695 -14.742 ;
      RECT 23.555 -15.515 23.695 -15.345 ;
      RECT 23.605 -14.328 23.695 -13.32 ;
      RECT 23.555 -13.725 23.695 -13.555 ;
      RECT 23.605 -12.52 23.695 -11.512 ;
      RECT 23.555 -12.285 23.695 -12.115 ;
      RECT 23.605 -11.098 23.695 -10.09 ;
      RECT 23.555 -10.495 23.695 -10.325 ;
      RECT 23.605 -9.29 23.695 -8.282 ;
      RECT 23.555 -9.055 23.695 -8.885 ;
      RECT 23.605 -7.868 23.695 -6.86 ;
      RECT 23.555 -7.265 23.695 -7.095 ;
      RECT 23.605 -6.06 23.695 -5.052 ;
      RECT 23.555 -5.825 23.695 -5.655 ;
      RECT 23.605 -4.638 23.695 -3.63 ;
      RECT 23.555 -4.035 23.695 -3.865 ;
      RECT 23.605 -2.83 23.695 -1.822 ;
      RECT 23.555 -2.595 23.695 -2.425 ;
      RECT 23.605 -1.408 23.695 -0.4 ;
      RECT 23.555 -0.805 23.695 -0.635 ;
      RECT 23.605 0.4 23.695 1.408 ;
      RECT 23.555 0.635 23.695 0.805 ;
      RECT 22.175 -60.005 23.655 -59.905 ;
      RECT 22.175 -60.515 22.275 -59.905 ;
      RECT 22.395 -57.47 23.655 -57.37 ;
      RECT 23.555 -57.795 23.655 -57.37 ;
      RECT 22.995 -57.795 23.095 -57.37 ;
      RECT 22.435 -57.795 22.535 -57.37 ;
      RECT 23.205 -49.858 23.295 -48.851 ;
      RECT 23.205 -49.545 23.345 -49.375 ;
      RECT 23.205 -48.049 23.295 -47.042 ;
      RECT 23.205 -47.525 23.345 -47.355 ;
      RECT 23.205 -46.628 23.295 -45.621 ;
      RECT 23.205 -46.315 23.345 -46.145 ;
      RECT 23.205 -44.819 23.295 -43.812 ;
      RECT 23.205 -44.295 23.345 -44.125 ;
      RECT 23.205 -43.398 23.295 -42.391 ;
      RECT 23.205 -43.085 23.345 -42.915 ;
      RECT 23.205 -41.589 23.295 -40.582 ;
      RECT 23.205 -41.065 23.345 -40.895 ;
      RECT 23.205 -40.168 23.295 -39.161 ;
      RECT 23.205 -39.855 23.345 -39.685 ;
      RECT 23.205 -38.359 23.295 -37.352 ;
      RECT 23.205 -37.835 23.345 -37.665 ;
      RECT 23.205 -36.938 23.295 -35.931 ;
      RECT 23.205 -36.625 23.345 -36.455 ;
      RECT 23.205 -35.129 23.295 -34.122 ;
      RECT 23.205 -34.605 23.345 -34.435 ;
      RECT 23.205 -33.708 23.295 -32.701 ;
      RECT 23.205 -33.395 23.345 -33.225 ;
      RECT 23.205 -31.899 23.295 -30.892 ;
      RECT 23.205 -31.375 23.345 -31.205 ;
      RECT 23.205 -30.478 23.295 -29.471 ;
      RECT 23.205 -30.165 23.345 -29.995 ;
      RECT 23.205 -28.669 23.295 -27.662 ;
      RECT 23.205 -28.145 23.345 -27.975 ;
      RECT 23.205 -27.248 23.295 -26.241 ;
      RECT 23.205 -26.935 23.345 -26.765 ;
      RECT 23.205 -25.439 23.295 -24.432 ;
      RECT 23.205 -24.915 23.345 -24.745 ;
      RECT 23.205 -24.018 23.295 -23.011 ;
      RECT 23.205 -23.705 23.345 -23.535 ;
      RECT 23.205 -22.209 23.295 -21.202 ;
      RECT 23.205 -21.685 23.345 -21.515 ;
      RECT 23.205 -20.788 23.295 -19.781 ;
      RECT 23.205 -20.475 23.345 -20.305 ;
      RECT 23.205 -18.979 23.295 -17.972 ;
      RECT 23.205 -18.455 23.345 -18.285 ;
      RECT 23.205 -17.558 23.295 -16.551 ;
      RECT 23.205 -17.245 23.345 -17.075 ;
      RECT 23.205 -15.749 23.295 -14.742 ;
      RECT 23.205 -15.225 23.345 -15.055 ;
      RECT 23.205 -14.328 23.295 -13.321 ;
      RECT 23.205 -14.015 23.345 -13.845 ;
      RECT 23.205 -12.519 23.295 -11.512 ;
      RECT 23.205 -11.995 23.345 -11.825 ;
      RECT 23.205 -11.098 23.295 -10.091 ;
      RECT 23.205 -10.785 23.345 -10.615 ;
      RECT 23.205 -9.289 23.295 -8.282 ;
      RECT 23.205 -8.765 23.345 -8.595 ;
      RECT 23.205 -7.868 23.295 -6.861 ;
      RECT 23.205 -7.555 23.345 -7.385 ;
      RECT 23.205 -6.059 23.295 -5.052 ;
      RECT 23.205 -5.535 23.345 -5.365 ;
      RECT 23.205 -4.638 23.295 -3.631 ;
      RECT 23.205 -4.325 23.345 -4.155 ;
      RECT 23.205 -2.829 23.295 -1.822 ;
      RECT 23.205 -2.305 23.345 -2.135 ;
      RECT 23.205 -1.408 23.295 -0.401 ;
      RECT 23.205 -1.095 23.345 -0.925 ;
      RECT 23.205 0.401 23.295 1.408 ;
      RECT 23.205 0.925 23.345 1.095 ;
      RECT 22.535 -59.815 22.705 -59.705 ;
      RECT 19.385 -59.815 22.705 -59.715 ;
      RECT 22.405 -49.858 22.495 -48.85 ;
      RECT 22.355 -49.255 22.495 -49.085 ;
      RECT 22.405 -48.05 22.495 -47.042 ;
      RECT 22.355 -47.815 22.495 -47.645 ;
      RECT 22.405 -46.628 22.495 -45.62 ;
      RECT 22.355 -46.025 22.495 -45.855 ;
      RECT 22.405 -44.82 22.495 -43.812 ;
      RECT 22.355 -44.585 22.495 -44.415 ;
      RECT 22.405 -43.398 22.495 -42.39 ;
      RECT 22.355 -42.795 22.495 -42.625 ;
      RECT 22.405 -41.59 22.495 -40.582 ;
      RECT 22.355 -41.355 22.495 -41.185 ;
      RECT 22.405 -40.168 22.495 -39.16 ;
      RECT 22.355 -39.565 22.495 -39.395 ;
      RECT 22.405 -38.36 22.495 -37.352 ;
      RECT 22.355 -38.125 22.495 -37.955 ;
      RECT 22.405 -36.938 22.495 -35.93 ;
      RECT 22.355 -36.335 22.495 -36.165 ;
      RECT 22.405 -35.13 22.495 -34.122 ;
      RECT 22.355 -34.895 22.495 -34.725 ;
      RECT 22.405 -33.708 22.495 -32.7 ;
      RECT 22.355 -33.105 22.495 -32.935 ;
      RECT 22.405 -31.9 22.495 -30.892 ;
      RECT 22.355 -31.665 22.495 -31.495 ;
      RECT 22.405 -30.478 22.495 -29.47 ;
      RECT 22.355 -29.875 22.495 -29.705 ;
      RECT 22.405 -28.67 22.495 -27.662 ;
      RECT 22.355 -28.435 22.495 -28.265 ;
      RECT 22.405 -27.248 22.495 -26.24 ;
      RECT 22.355 -26.645 22.495 -26.475 ;
      RECT 22.405 -25.44 22.495 -24.432 ;
      RECT 22.355 -25.205 22.495 -25.035 ;
      RECT 22.405 -24.018 22.495 -23.01 ;
      RECT 22.355 -23.415 22.495 -23.245 ;
      RECT 22.405 -22.21 22.495 -21.202 ;
      RECT 22.355 -21.975 22.495 -21.805 ;
      RECT 22.405 -20.788 22.495 -19.78 ;
      RECT 22.355 -20.185 22.495 -20.015 ;
      RECT 22.405 -18.98 22.495 -17.972 ;
      RECT 22.355 -18.745 22.495 -18.575 ;
      RECT 22.405 -17.558 22.495 -16.55 ;
      RECT 22.355 -16.955 22.495 -16.785 ;
      RECT 22.405 -15.75 22.495 -14.742 ;
      RECT 22.355 -15.515 22.495 -15.345 ;
      RECT 22.405 -14.328 22.495 -13.32 ;
      RECT 22.355 -13.725 22.495 -13.555 ;
      RECT 22.405 -12.52 22.495 -11.512 ;
      RECT 22.355 -12.285 22.495 -12.115 ;
      RECT 22.405 -11.098 22.495 -10.09 ;
      RECT 22.355 -10.495 22.495 -10.325 ;
      RECT 22.405 -9.29 22.495 -8.282 ;
      RECT 22.355 -9.055 22.495 -8.885 ;
      RECT 22.405 -7.868 22.495 -6.86 ;
      RECT 22.355 -7.265 22.495 -7.095 ;
      RECT 22.405 -6.06 22.495 -5.052 ;
      RECT 22.355 -5.825 22.495 -5.655 ;
      RECT 22.405 -4.638 22.495 -3.63 ;
      RECT 22.355 -4.035 22.495 -3.865 ;
      RECT 22.405 -2.83 22.495 -1.822 ;
      RECT 22.355 -2.595 22.495 -2.425 ;
      RECT 22.405 -1.408 22.495 -0.4 ;
      RECT 22.355 -0.805 22.495 -0.635 ;
      RECT 22.405 0.4 22.495 1.408 ;
      RECT 22.355 0.635 22.495 0.805 ;
      RECT 22.005 -49.858 22.095 -48.851 ;
      RECT 22.005 -49.545 22.145 -49.375 ;
      RECT 22.005 -48.049 22.095 -47.042 ;
      RECT 22.005 -47.525 22.145 -47.355 ;
      RECT 22.005 -46.628 22.095 -45.621 ;
      RECT 22.005 -46.315 22.145 -46.145 ;
      RECT 22.005 -44.819 22.095 -43.812 ;
      RECT 22.005 -44.295 22.145 -44.125 ;
      RECT 22.005 -43.398 22.095 -42.391 ;
      RECT 22.005 -43.085 22.145 -42.915 ;
      RECT 22.005 -41.589 22.095 -40.582 ;
      RECT 22.005 -41.065 22.145 -40.895 ;
      RECT 22.005 -40.168 22.095 -39.161 ;
      RECT 22.005 -39.855 22.145 -39.685 ;
      RECT 22.005 -38.359 22.095 -37.352 ;
      RECT 22.005 -37.835 22.145 -37.665 ;
      RECT 22.005 -36.938 22.095 -35.931 ;
      RECT 22.005 -36.625 22.145 -36.455 ;
      RECT 22.005 -35.129 22.095 -34.122 ;
      RECT 22.005 -34.605 22.145 -34.435 ;
      RECT 22.005 -33.708 22.095 -32.701 ;
      RECT 22.005 -33.395 22.145 -33.225 ;
      RECT 22.005 -31.899 22.095 -30.892 ;
      RECT 22.005 -31.375 22.145 -31.205 ;
      RECT 22.005 -30.478 22.095 -29.471 ;
      RECT 22.005 -30.165 22.145 -29.995 ;
      RECT 22.005 -28.669 22.095 -27.662 ;
      RECT 22.005 -28.145 22.145 -27.975 ;
      RECT 22.005 -27.248 22.095 -26.241 ;
      RECT 22.005 -26.935 22.145 -26.765 ;
      RECT 22.005 -25.439 22.095 -24.432 ;
      RECT 22.005 -24.915 22.145 -24.745 ;
      RECT 22.005 -24.018 22.095 -23.011 ;
      RECT 22.005 -23.705 22.145 -23.535 ;
      RECT 22.005 -22.209 22.095 -21.202 ;
      RECT 22.005 -21.685 22.145 -21.515 ;
      RECT 22.005 -20.788 22.095 -19.781 ;
      RECT 22.005 -20.475 22.145 -20.305 ;
      RECT 22.005 -18.979 22.095 -17.972 ;
      RECT 22.005 -18.455 22.145 -18.285 ;
      RECT 22.005 -17.558 22.095 -16.551 ;
      RECT 22.005 -17.245 22.145 -17.075 ;
      RECT 22.005 -15.749 22.095 -14.742 ;
      RECT 22.005 -15.225 22.145 -15.055 ;
      RECT 22.005 -14.328 22.095 -13.321 ;
      RECT 22.005 -14.015 22.145 -13.845 ;
      RECT 22.005 -12.519 22.095 -11.512 ;
      RECT 22.005 -11.995 22.145 -11.825 ;
      RECT 22.005 -11.098 22.095 -10.091 ;
      RECT 22.005 -10.785 22.145 -10.615 ;
      RECT 22.005 -9.289 22.095 -8.282 ;
      RECT 22.005 -8.765 22.145 -8.595 ;
      RECT 22.005 -7.868 22.095 -6.861 ;
      RECT 22.005 -7.555 22.145 -7.385 ;
      RECT 22.005 -6.059 22.095 -5.052 ;
      RECT 22.005 -5.535 22.145 -5.365 ;
      RECT 22.005 -4.638 22.095 -3.631 ;
      RECT 22.005 -4.325 22.145 -4.155 ;
      RECT 22.005 -2.829 22.095 -1.822 ;
      RECT 22.005 -2.305 22.145 -2.135 ;
      RECT 22.005 -1.408 22.095 -0.401 ;
      RECT 22.005 -1.095 22.145 -0.925 ;
      RECT 22.005 0.401 22.095 1.408 ;
      RECT 22.005 0.925 22.145 1.095 ;
      RECT 20.155 -60.005 21.635 -59.905 ;
      RECT 20.155 -60.375 20.255 -59.905 ;
      RECT 19.96 -62.715 21.535 -62.595 ;
      RECT 21.435 -63.215 21.535 -62.595 ;
      RECT 20.84 -63.215 20.94 -62.595 ;
      RECT 19.96 -63.17 20.06 -62.595 ;
      RECT 21.205 -49.858 21.295 -48.85 ;
      RECT 21.155 -49.255 21.295 -49.085 ;
      RECT 21.205 -48.05 21.295 -47.042 ;
      RECT 21.155 -47.815 21.295 -47.645 ;
      RECT 21.205 -46.628 21.295 -45.62 ;
      RECT 21.155 -46.025 21.295 -45.855 ;
      RECT 21.205 -44.82 21.295 -43.812 ;
      RECT 21.155 -44.585 21.295 -44.415 ;
      RECT 21.205 -43.398 21.295 -42.39 ;
      RECT 21.155 -42.795 21.295 -42.625 ;
      RECT 21.205 -41.59 21.295 -40.582 ;
      RECT 21.155 -41.355 21.295 -41.185 ;
      RECT 21.205 -40.168 21.295 -39.16 ;
      RECT 21.155 -39.565 21.295 -39.395 ;
      RECT 21.205 -38.36 21.295 -37.352 ;
      RECT 21.155 -38.125 21.295 -37.955 ;
      RECT 21.205 -36.938 21.295 -35.93 ;
      RECT 21.155 -36.335 21.295 -36.165 ;
      RECT 21.205 -35.13 21.295 -34.122 ;
      RECT 21.155 -34.895 21.295 -34.725 ;
      RECT 21.205 -33.708 21.295 -32.7 ;
      RECT 21.155 -33.105 21.295 -32.935 ;
      RECT 21.205 -31.9 21.295 -30.892 ;
      RECT 21.155 -31.665 21.295 -31.495 ;
      RECT 21.205 -30.478 21.295 -29.47 ;
      RECT 21.155 -29.875 21.295 -29.705 ;
      RECT 21.205 -28.67 21.295 -27.662 ;
      RECT 21.155 -28.435 21.295 -28.265 ;
      RECT 21.205 -27.248 21.295 -26.24 ;
      RECT 21.155 -26.645 21.295 -26.475 ;
      RECT 21.205 -25.44 21.295 -24.432 ;
      RECT 21.155 -25.205 21.295 -25.035 ;
      RECT 21.205 -24.018 21.295 -23.01 ;
      RECT 21.155 -23.415 21.295 -23.245 ;
      RECT 21.205 -22.21 21.295 -21.202 ;
      RECT 21.155 -21.975 21.295 -21.805 ;
      RECT 21.205 -20.788 21.295 -19.78 ;
      RECT 21.155 -20.185 21.295 -20.015 ;
      RECT 21.205 -18.98 21.295 -17.972 ;
      RECT 21.155 -18.745 21.295 -18.575 ;
      RECT 21.205 -17.558 21.295 -16.55 ;
      RECT 21.155 -16.955 21.295 -16.785 ;
      RECT 21.205 -15.75 21.295 -14.742 ;
      RECT 21.155 -15.515 21.295 -15.345 ;
      RECT 21.205 -14.328 21.295 -13.32 ;
      RECT 21.155 -13.725 21.295 -13.555 ;
      RECT 21.205 -12.52 21.295 -11.512 ;
      RECT 21.155 -12.285 21.295 -12.115 ;
      RECT 21.205 -11.098 21.295 -10.09 ;
      RECT 21.155 -10.495 21.295 -10.325 ;
      RECT 21.205 -9.29 21.295 -8.282 ;
      RECT 21.155 -9.055 21.295 -8.885 ;
      RECT 21.205 -7.868 21.295 -6.86 ;
      RECT 21.155 -7.265 21.295 -7.095 ;
      RECT 21.205 -6.06 21.295 -5.052 ;
      RECT 21.155 -5.825 21.295 -5.655 ;
      RECT 21.205 -4.638 21.295 -3.63 ;
      RECT 21.155 -4.035 21.295 -3.865 ;
      RECT 21.205 -2.83 21.295 -1.822 ;
      RECT 21.155 -2.595 21.295 -2.425 ;
      RECT 21.205 -1.408 21.295 -0.4 ;
      RECT 21.155 -0.805 21.295 -0.635 ;
      RECT 21.205 0.4 21.295 1.408 ;
      RECT 21.155 0.635 21.295 0.805 ;
      RECT 21.08 -63.005 21.255 -62.835 ;
      RECT 21.155 -63.215 21.255 -62.835 ;
      RECT 20.195 -61.875 20.295 -61.41 ;
      RECT 20.56 -61.875 20.66 -61.42 ;
      RECT 20.195 -61.875 21.04 -61.705 ;
      RECT 20.805 -49.858 20.895 -48.851 ;
      RECT 20.805 -49.545 20.945 -49.375 ;
      RECT 20.805 -48.049 20.895 -47.042 ;
      RECT 20.805 -47.525 20.945 -47.355 ;
      RECT 20.805 -46.628 20.895 -45.621 ;
      RECT 20.805 -46.315 20.945 -46.145 ;
      RECT 20.805 -44.819 20.895 -43.812 ;
      RECT 20.805 -44.295 20.945 -44.125 ;
      RECT 20.805 -43.398 20.895 -42.391 ;
      RECT 20.805 -43.085 20.945 -42.915 ;
      RECT 20.805 -41.589 20.895 -40.582 ;
      RECT 20.805 -41.065 20.945 -40.895 ;
      RECT 20.805 -40.168 20.895 -39.161 ;
      RECT 20.805 -39.855 20.945 -39.685 ;
      RECT 20.805 -38.359 20.895 -37.352 ;
      RECT 20.805 -37.835 20.945 -37.665 ;
      RECT 20.805 -36.938 20.895 -35.931 ;
      RECT 20.805 -36.625 20.945 -36.455 ;
      RECT 20.805 -35.129 20.895 -34.122 ;
      RECT 20.805 -34.605 20.945 -34.435 ;
      RECT 20.805 -33.708 20.895 -32.701 ;
      RECT 20.805 -33.395 20.945 -33.225 ;
      RECT 20.805 -31.899 20.895 -30.892 ;
      RECT 20.805 -31.375 20.945 -31.205 ;
      RECT 20.805 -30.478 20.895 -29.471 ;
      RECT 20.805 -30.165 20.945 -29.995 ;
      RECT 20.805 -28.669 20.895 -27.662 ;
      RECT 20.805 -28.145 20.945 -27.975 ;
      RECT 20.805 -27.248 20.895 -26.241 ;
      RECT 20.805 -26.935 20.945 -26.765 ;
      RECT 20.805 -25.439 20.895 -24.432 ;
      RECT 20.805 -24.915 20.945 -24.745 ;
      RECT 20.805 -24.018 20.895 -23.011 ;
      RECT 20.805 -23.705 20.945 -23.535 ;
      RECT 20.805 -22.209 20.895 -21.202 ;
      RECT 20.805 -21.685 20.945 -21.515 ;
      RECT 20.805 -20.788 20.895 -19.781 ;
      RECT 20.805 -20.475 20.945 -20.305 ;
      RECT 20.805 -18.979 20.895 -17.972 ;
      RECT 20.805 -18.455 20.945 -18.285 ;
      RECT 20.805 -17.558 20.895 -16.551 ;
      RECT 20.805 -17.245 20.945 -17.075 ;
      RECT 20.805 -15.749 20.895 -14.742 ;
      RECT 20.805 -15.225 20.945 -15.055 ;
      RECT 20.805 -14.328 20.895 -13.321 ;
      RECT 20.805 -14.015 20.945 -13.845 ;
      RECT 20.805 -12.519 20.895 -11.512 ;
      RECT 20.805 -11.995 20.945 -11.825 ;
      RECT 20.805 -11.098 20.895 -10.091 ;
      RECT 20.805 -10.785 20.945 -10.615 ;
      RECT 20.805 -9.289 20.895 -8.282 ;
      RECT 20.805 -8.765 20.945 -8.595 ;
      RECT 20.805 -7.868 20.895 -6.861 ;
      RECT 20.805 -7.555 20.945 -7.385 ;
      RECT 20.805 -6.059 20.895 -5.052 ;
      RECT 20.805 -5.535 20.945 -5.365 ;
      RECT 20.805 -4.638 20.895 -3.631 ;
      RECT 20.805 -4.325 20.945 -4.155 ;
      RECT 20.805 -2.829 20.895 -1.822 ;
      RECT 20.805 -2.305 20.945 -2.135 ;
      RECT 20.805 -1.408 20.895 -0.401 ;
      RECT 20.805 -1.095 20.945 -0.925 ;
      RECT 20.805 0.401 20.895 1.408 ;
      RECT 20.805 0.925 20.945 1.095 ;
      RECT 20.49 -63.005 20.66 -62.835 ;
      RECT 20.56 -63.215 20.66 -62.835 ;
      RECT 20.005 -49.858 20.095 -48.85 ;
      RECT 19.955 -49.255 20.095 -49.085 ;
      RECT 20.005 -48.05 20.095 -47.042 ;
      RECT 19.955 -47.815 20.095 -47.645 ;
      RECT 20.005 -46.628 20.095 -45.62 ;
      RECT 19.955 -46.025 20.095 -45.855 ;
      RECT 20.005 -44.82 20.095 -43.812 ;
      RECT 19.955 -44.585 20.095 -44.415 ;
      RECT 20.005 -43.398 20.095 -42.39 ;
      RECT 19.955 -42.795 20.095 -42.625 ;
      RECT 20.005 -41.59 20.095 -40.582 ;
      RECT 19.955 -41.355 20.095 -41.185 ;
      RECT 20.005 -40.168 20.095 -39.16 ;
      RECT 19.955 -39.565 20.095 -39.395 ;
      RECT 20.005 -38.36 20.095 -37.352 ;
      RECT 19.955 -38.125 20.095 -37.955 ;
      RECT 20.005 -36.938 20.095 -35.93 ;
      RECT 19.955 -36.335 20.095 -36.165 ;
      RECT 20.005 -35.13 20.095 -34.122 ;
      RECT 19.955 -34.895 20.095 -34.725 ;
      RECT 20.005 -33.708 20.095 -32.7 ;
      RECT 19.955 -33.105 20.095 -32.935 ;
      RECT 20.005 -31.9 20.095 -30.892 ;
      RECT 19.955 -31.665 20.095 -31.495 ;
      RECT 20.005 -30.478 20.095 -29.47 ;
      RECT 19.955 -29.875 20.095 -29.705 ;
      RECT 20.005 -28.67 20.095 -27.662 ;
      RECT 19.955 -28.435 20.095 -28.265 ;
      RECT 20.005 -27.248 20.095 -26.24 ;
      RECT 19.955 -26.645 20.095 -26.475 ;
      RECT 20.005 -25.44 20.095 -24.432 ;
      RECT 19.955 -25.205 20.095 -25.035 ;
      RECT 20.005 -24.018 20.095 -23.01 ;
      RECT 19.955 -23.415 20.095 -23.245 ;
      RECT 20.005 -22.21 20.095 -21.202 ;
      RECT 19.955 -21.975 20.095 -21.805 ;
      RECT 20.005 -20.788 20.095 -19.78 ;
      RECT 19.955 -20.185 20.095 -20.015 ;
      RECT 20.005 -18.98 20.095 -17.972 ;
      RECT 19.955 -18.745 20.095 -18.575 ;
      RECT 20.005 -17.558 20.095 -16.55 ;
      RECT 19.955 -16.955 20.095 -16.785 ;
      RECT 20.005 -15.75 20.095 -14.742 ;
      RECT 19.955 -15.515 20.095 -15.345 ;
      RECT 20.005 -14.328 20.095 -13.32 ;
      RECT 19.955 -13.725 20.095 -13.555 ;
      RECT 20.005 -12.52 20.095 -11.512 ;
      RECT 19.955 -12.285 20.095 -12.115 ;
      RECT 20.005 -11.098 20.095 -10.09 ;
      RECT 19.955 -10.495 20.095 -10.325 ;
      RECT 20.005 -9.29 20.095 -8.282 ;
      RECT 19.955 -9.055 20.095 -8.885 ;
      RECT 20.005 -7.868 20.095 -6.86 ;
      RECT 19.955 -7.265 20.095 -7.095 ;
      RECT 20.005 -6.06 20.095 -5.052 ;
      RECT 19.955 -5.825 20.095 -5.655 ;
      RECT 20.005 -4.638 20.095 -3.63 ;
      RECT 19.955 -4.035 20.095 -3.865 ;
      RECT 20.005 -2.83 20.095 -1.822 ;
      RECT 19.955 -2.595 20.095 -2.425 ;
      RECT 20.005 -1.408 20.095 -0.4 ;
      RECT 19.955 -0.805 20.095 -0.635 ;
      RECT 20.005 0.4 20.095 1.408 ;
      RECT 19.955 0.635 20.095 0.805 ;
      RECT 19.605 -49.858 19.695 -48.851 ;
      RECT 19.605 -49.545 19.745 -49.375 ;
      RECT 19.605 -48.049 19.695 -47.042 ;
      RECT 19.605 -47.525 19.745 -47.355 ;
      RECT 19.605 -46.628 19.695 -45.621 ;
      RECT 19.605 -46.315 19.745 -46.145 ;
      RECT 19.605 -44.819 19.695 -43.812 ;
      RECT 19.605 -44.295 19.745 -44.125 ;
      RECT 19.605 -43.398 19.695 -42.391 ;
      RECT 19.605 -43.085 19.745 -42.915 ;
      RECT 19.605 -41.589 19.695 -40.582 ;
      RECT 19.605 -41.065 19.745 -40.895 ;
      RECT 19.605 -40.168 19.695 -39.161 ;
      RECT 19.605 -39.855 19.745 -39.685 ;
      RECT 19.605 -38.359 19.695 -37.352 ;
      RECT 19.605 -37.835 19.745 -37.665 ;
      RECT 19.605 -36.938 19.695 -35.931 ;
      RECT 19.605 -36.625 19.745 -36.455 ;
      RECT 19.605 -35.129 19.695 -34.122 ;
      RECT 19.605 -34.605 19.745 -34.435 ;
      RECT 19.605 -33.708 19.695 -32.701 ;
      RECT 19.605 -33.395 19.745 -33.225 ;
      RECT 19.605 -31.899 19.695 -30.892 ;
      RECT 19.605 -31.375 19.745 -31.205 ;
      RECT 19.605 -30.478 19.695 -29.471 ;
      RECT 19.605 -30.165 19.745 -29.995 ;
      RECT 19.605 -28.669 19.695 -27.662 ;
      RECT 19.605 -28.145 19.745 -27.975 ;
      RECT 19.605 -27.248 19.695 -26.241 ;
      RECT 19.605 -26.935 19.745 -26.765 ;
      RECT 19.605 -25.439 19.695 -24.432 ;
      RECT 19.605 -24.915 19.745 -24.745 ;
      RECT 19.605 -24.018 19.695 -23.011 ;
      RECT 19.605 -23.705 19.745 -23.535 ;
      RECT 19.605 -22.209 19.695 -21.202 ;
      RECT 19.605 -21.685 19.745 -21.515 ;
      RECT 19.605 -20.788 19.695 -19.781 ;
      RECT 19.605 -20.475 19.745 -20.305 ;
      RECT 19.605 -18.979 19.695 -17.972 ;
      RECT 19.605 -18.455 19.745 -18.285 ;
      RECT 19.605 -17.558 19.695 -16.551 ;
      RECT 19.605 -17.245 19.745 -17.075 ;
      RECT 19.605 -15.749 19.695 -14.742 ;
      RECT 19.605 -15.225 19.745 -15.055 ;
      RECT 19.605 -14.328 19.695 -13.321 ;
      RECT 19.605 -14.015 19.745 -13.845 ;
      RECT 19.605 -12.519 19.695 -11.512 ;
      RECT 19.605 -11.995 19.745 -11.825 ;
      RECT 19.605 -11.098 19.695 -10.091 ;
      RECT 19.605 -10.785 19.745 -10.615 ;
      RECT 19.605 -9.289 19.695 -8.282 ;
      RECT 19.605 -8.765 19.745 -8.595 ;
      RECT 19.605 -7.868 19.695 -6.861 ;
      RECT 19.605 -7.555 19.745 -7.385 ;
      RECT 19.605 -6.059 19.695 -5.052 ;
      RECT 19.605 -5.535 19.745 -5.365 ;
      RECT 19.605 -4.638 19.695 -3.631 ;
      RECT 19.605 -4.325 19.745 -4.155 ;
      RECT 19.605 -2.829 19.695 -1.822 ;
      RECT 19.605 -2.305 19.745 -2.135 ;
      RECT 19.605 -1.408 19.695 -0.401 ;
      RECT 19.605 -1.095 19.745 -0.925 ;
      RECT 19.605 0.401 19.695 1.408 ;
      RECT 19.605 0.925 19.745 1.095 ;
      RECT 15.435 -57.255 19.215 -57.135 ;
      RECT 16.755 -57.795 16.855 -57.135 ;
      RECT 16.195 -57.795 16.295 -57.135 ;
      RECT 15.635 -57.795 15.735 -57.135 ;
      RECT 18.805 -49.858 18.895 -48.85 ;
      RECT 18.755 -49.255 18.895 -49.085 ;
      RECT 18.805 -48.05 18.895 -47.042 ;
      RECT 18.755 -47.815 18.895 -47.645 ;
      RECT 18.805 -46.628 18.895 -45.62 ;
      RECT 18.755 -46.025 18.895 -45.855 ;
      RECT 18.805 -44.82 18.895 -43.812 ;
      RECT 18.755 -44.585 18.895 -44.415 ;
      RECT 18.805 -43.398 18.895 -42.39 ;
      RECT 18.755 -42.795 18.895 -42.625 ;
      RECT 18.805 -41.59 18.895 -40.582 ;
      RECT 18.755 -41.355 18.895 -41.185 ;
      RECT 18.805 -40.168 18.895 -39.16 ;
      RECT 18.755 -39.565 18.895 -39.395 ;
      RECT 18.805 -38.36 18.895 -37.352 ;
      RECT 18.755 -38.125 18.895 -37.955 ;
      RECT 18.805 -36.938 18.895 -35.93 ;
      RECT 18.755 -36.335 18.895 -36.165 ;
      RECT 18.805 -35.13 18.895 -34.122 ;
      RECT 18.755 -34.895 18.895 -34.725 ;
      RECT 18.805 -33.708 18.895 -32.7 ;
      RECT 18.755 -33.105 18.895 -32.935 ;
      RECT 18.805 -31.9 18.895 -30.892 ;
      RECT 18.755 -31.665 18.895 -31.495 ;
      RECT 18.805 -30.478 18.895 -29.47 ;
      RECT 18.755 -29.875 18.895 -29.705 ;
      RECT 18.805 -28.67 18.895 -27.662 ;
      RECT 18.755 -28.435 18.895 -28.265 ;
      RECT 18.805 -27.248 18.895 -26.24 ;
      RECT 18.755 -26.645 18.895 -26.475 ;
      RECT 18.805 -25.44 18.895 -24.432 ;
      RECT 18.755 -25.205 18.895 -25.035 ;
      RECT 18.805 -24.018 18.895 -23.01 ;
      RECT 18.755 -23.415 18.895 -23.245 ;
      RECT 18.805 -22.21 18.895 -21.202 ;
      RECT 18.755 -21.975 18.895 -21.805 ;
      RECT 18.805 -20.788 18.895 -19.78 ;
      RECT 18.755 -20.185 18.895 -20.015 ;
      RECT 18.805 -18.98 18.895 -17.972 ;
      RECT 18.755 -18.745 18.895 -18.575 ;
      RECT 18.805 -17.558 18.895 -16.55 ;
      RECT 18.755 -16.955 18.895 -16.785 ;
      RECT 18.805 -15.75 18.895 -14.742 ;
      RECT 18.755 -15.515 18.895 -15.345 ;
      RECT 18.805 -14.328 18.895 -13.32 ;
      RECT 18.755 -13.725 18.895 -13.555 ;
      RECT 18.805 -12.52 18.895 -11.512 ;
      RECT 18.755 -12.285 18.895 -12.115 ;
      RECT 18.805 -11.098 18.895 -10.09 ;
      RECT 18.755 -10.495 18.895 -10.325 ;
      RECT 18.805 -9.29 18.895 -8.282 ;
      RECT 18.755 -9.055 18.895 -8.885 ;
      RECT 18.805 -7.868 18.895 -6.86 ;
      RECT 18.755 -7.265 18.895 -7.095 ;
      RECT 18.805 -6.06 18.895 -5.052 ;
      RECT 18.755 -5.825 18.895 -5.655 ;
      RECT 18.805 -4.638 18.895 -3.63 ;
      RECT 18.755 -4.035 18.895 -3.865 ;
      RECT 18.805 -2.83 18.895 -1.822 ;
      RECT 18.755 -2.595 18.895 -2.425 ;
      RECT 18.805 -1.408 18.895 -0.4 ;
      RECT 18.755 -0.805 18.895 -0.635 ;
      RECT 18.805 0.4 18.895 1.408 ;
      RECT 18.755 0.635 18.895 0.805 ;
      RECT 17.375 -60.005 18.855 -59.905 ;
      RECT 17.375 -60.515 17.475 -59.905 ;
      RECT 17.595 -57.47 18.855 -57.37 ;
      RECT 18.755 -57.795 18.855 -57.37 ;
      RECT 18.195 -57.795 18.295 -57.37 ;
      RECT 17.635 -57.795 17.735 -57.37 ;
      RECT 18.405 -49.858 18.495 -48.851 ;
      RECT 18.405 -49.545 18.545 -49.375 ;
      RECT 18.405 -48.049 18.495 -47.042 ;
      RECT 18.405 -47.525 18.545 -47.355 ;
      RECT 18.405 -46.628 18.495 -45.621 ;
      RECT 18.405 -46.315 18.545 -46.145 ;
      RECT 18.405 -44.819 18.495 -43.812 ;
      RECT 18.405 -44.295 18.545 -44.125 ;
      RECT 18.405 -43.398 18.495 -42.391 ;
      RECT 18.405 -43.085 18.545 -42.915 ;
      RECT 18.405 -41.589 18.495 -40.582 ;
      RECT 18.405 -41.065 18.545 -40.895 ;
      RECT 18.405 -40.168 18.495 -39.161 ;
      RECT 18.405 -39.855 18.545 -39.685 ;
      RECT 18.405 -38.359 18.495 -37.352 ;
      RECT 18.405 -37.835 18.545 -37.665 ;
      RECT 18.405 -36.938 18.495 -35.931 ;
      RECT 18.405 -36.625 18.545 -36.455 ;
      RECT 18.405 -35.129 18.495 -34.122 ;
      RECT 18.405 -34.605 18.545 -34.435 ;
      RECT 18.405 -33.708 18.495 -32.701 ;
      RECT 18.405 -33.395 18.545 -33.225 ;
      RECT 18.405 -31.899 18.495 -30.892 ;
      RECT 18.405 -31.375 18.545 -31.205 ;
      RECT 18.405 -30.478 18.495 -29.471 ;
      RECT 18.405 -30.165 18.545 -29.995 ;
      RECT 18.405 -28.669 18.495 -27.662 ;
      RECT 18.405 -28.145 18.545 -27.975 ;
      RECT 18.405 -27.248 18.495 -26.241 ;
      RECT 18.405 -26.935 18.545 -26.765 ;
      RECT 18.405 -25.439 18.495 -24.432 ;
      RECT 18.405 -24.915 18.545 -24.745 ;
      RECT 18.405 -24.018 18.495 -23.011 ;
      RECT 18.405 -23.705 18.545 -23.535 ;
      RECT 18.405 -22.209 18.495 -21.202 ;
      RECT 18.405 -21.685 18.545 -21.515 ;
      RECT 18.405 -20.788 18.495 -19.781 ;
      RECT 18.405 -20.475 18.545 -20.305 ;
      RECT 18.405 -18.979 18.495 -17.972 ;
      RECT 18.405 -18.455 18.545 -18.285 ;
      RECT 18.405 -17.558 18.495 -16.551 ;
      RECT 18.405 -17.245 18.545 -17.075 ;
      RECT 18.405 -15.749 18.495 -14.742 ;
      RECT 18.405 -15.225 18.545 -15.055 ;
      RECT 18.405 -14.328 18.495 -13.321 ;
      RECT 18.405 -14.015 18.545 -13.845 ;
      RECT 18.405 -12.519 18.495 -11.512 ;
      RECT 18.405 -11.995 18.545 -11.825 ;
      RECT 18.405 -11.098 18.495 -10.091 ;
      RECT 18.405 -10.785 18.545 -10.615 ;
      RECT 18.405 -9.289 18.495 -8.282 ;
      RECT 18.405 -8.765 18.545 -8.595 ;
      RECT 18.405 -7.868 18.495 -6.861 ;
      RECT 18.405 -7.555 18.545 -7.385 ;
      RECT 18.405 -6.059 18.495 -5.052 ;
      RECT 18.405 -5.535 18.545 -5.365 ;
      RECT 18.405 -4.638 18.495 -3.631 ;
      RECT 18.405 -4.325 18.545 -4.155 ;
      RECT 18.405 -2.829 18.495 -1.822 ;
      RECT 18.405 -2.305 18.545 -2.135 ;
      RECT 18.405 -1.408 18.495 -0.401 ;
      RECT 18.405 -1.095 18.545 -0.925 ;
      RECT 18.405 0.401 18.495 1.408 ;
      RECT 18.405 0.925 18.545 1.095 ;
      RECT 17.735 -59.815 17.905 -59.705 ;
      RECT 14.585 -59.815 17.905 -59.715 ;
      RECT 17.605 -49.858 17.695 -48.85 ;
      RECT 17.555 -49.255 17.695 -49.085 ;
      RECT 17.605 -48.05 17.695 -47.042 ;
      RECT 17.555 -47.815 17.695 -47.645 ;
      RECT 17.605 -46.628 17.695 -45.62 ;
      RECT 17.555 -46.025 17.695 -45.855 ;
      RECT 17.605 -44.82 17.695 -43.812 ;
      RECT 17.555 -44.585 17.695 -44.415 ;
      RECT 17.605 -43.398 17.695 -42.39 ;
      RECT 17.555 -42.795 17.695 -42.625 ;
      RECT 17.605 -41.59 17.695 -40.582 ;
      RECT 17.555 -41.355 17.695 -41.185 ;
      RECT 17.605 -40.168 17.695 -39.16 ;
      RECT 17.555 -39.565 17.695 -39.395 ;
      RECT 17.605 -38.36 17.695 -37.352 ;
      RECT 17.555 -38.125 17.695 -37.955 ;
      RECT 17.605 -36.938 17.695 -35.93 ;
      RECT 17.555 -36.335 17.695 -36.165 ;
      RECT 17.605 -35.13 17.695 -34.122 ;
      RECT 17.555 -34.895 17.695 -34.725 ;
      RECT 17.605 -33.708 17.695 -32.7 ;
      RECT 17.555 -33.105 17.695 -32.935 ;
      RECT 17.605 -31.9 17.695 -30.892 ;
      RECT 17.555 -31.665 17.695 -31.495 ;
      RECT 17.605 -30.478 17.695 -29.47 ;
      RECT 17.555 -29.875 17.695 -29.705 ;
      RECT 17.605 -28.67 17.695 -27.662 ;
      RECT 17.555 -28.435 17.695 -28.265 ;
      RECT 17.605 -27.248 17.695 -26.24 ;
      RECT 17.555 -26.645 17.695 -26.475 ;
      RECT 17.605 -25.44 17.695 -24.432 ;
      RECT 17.555 -25.205 17.695 -25.035 ;
      RECT 17.605 -24.018 17.695 -23.01 ;
      RECT 17.555 -23.415 17.695 -23.245 ;
      RECT 17.605 -22.21 17.695 -21.202 ;
      RECT 17.555 -21.975 17.695 -21.805 ;
      RECT 17.605 -20.788 17.695 -19.78 ;
      RECT 17.555 -20.185 17.695 -20.015 ;
      RECT 17.605 -18.98 17.695 -17.972 ;
      RECT 17.555 -18.745 17.695 -18.575 ;
      RECT 17.605 -17.558 17.695 -16.55 ;
      RECT 17.555 -16.955 17.695 -16.785 ;
      RECT 17.605 -15.75 17.695 -14.742 ;
      RECT 17.555 -15.515 17.695 -15.345 ;
      RECT 17.605 -14.328 17.695 -13.32 ;
      RECT 17.555 -13.725 17.695 -13.555 ;
      RECT 17.605 -12.52 17.695 -11.512 ;
      RECT 17.555 -12.285 17.695 -12.115 ;
      RECT 17.605 -11.098 17.695 -10.09 ;
      RECT 17.555 -10.495 17.695 -10.325 ;
      RECT 17.605 -9.29 17.695 -8.282 ;
      RECT 17.555 -9.055 17.695 -8.885 ;
      RECT 17.605 -7.868 17.695 -6.86 ;
      RECT 17.555 -7.265 17.695 -7.095 ;
      RECT 17.605 -6.06 17.695 -5.052 ;
      RECT 17.555 -5.825 17.695 -5.655 ;
      RECT 17.605 -4.638 17.695 -3.63 ;
      RECT 17.555 -4.035 17.695 -3.865 ;
      RECT 17.605 -2.83 17.695 -1.822 ;
      RECT 17.555 -2.595 17.695 -2.425 ;
      RECT 17.605 -1.408 17.695 -0.4 ;
      RECT 17.555 -0.805 17.695 -0.635 ;
      RECT 17.605 0.4 17.695 1.408 ;
      RECT 17.555 0.635 17.695 0.805 ;
      RECT 17.205 -49.858 17.295 -48.851 ;
      RECT 17.205 -49.545 17.345 -49.375 ;
      RECT 17.205 -48.049 17.295 -47.042 ;
      RECT 17.205 -47.525 17.345 -47.355 ;
      RECT 17.205 -46.628 17.295 -45.621 ;
      RECT 17.205 -46.315 17.345 -46.145 ;
      RECT 17.205 -44.819 17.295 -43.812 ;
      RECT 17.205 -44.295 17.345 -44.125 ;
      RECT 17.205 -43.398 17.295 -42.391 ;
      RECT 17.205 -43.085 17.345 -42.915 ;
      RECT 17.205 -41.589 17.295 -40.582 ;
      RECT 17.205 -41.065 17.345 -40.895 ;
      RECT 17.205 -40.168 17.295 -39.161 ;
      RECT 17.205 -39.855 17.345 -39.685 ;
      RECT 17.205 -38.359 17.295 -37.352 ;
      RECT 17.205 -37.835 17.345 -37.665 ;
      RECT 17.205 -36.938 17.295 -35.931 ;
      RECT 17.205 -36.625 17.345 -36.455 ;
      RECT 17.205 -35.129 17.295 -34.122 ;
      RECT 17.205 -34.605 17.345 -34.435 ;
      RECT 17.205 -33.708 17.295 -32.701 ;
      RECT 17.205 -33.395 17.345 -33.225 ;
      RECT 17.205 -31.899 17.295 -30.892 ;
      RECT 17.205 -31.375 17.345 -31.205 ;
      RECT 17.205 -30.478 17.295 -29.471 ;
      RECT 17.205 -30.165 17.345 -29.995 ;
      RECT 17.205 -28.669 17.295 -27.662 ;
      RECT 17.205 -28.145 17.345 -27.975 ;
      RECT 17.205 -27.248 17.295 -26.241 ;
      RECT 17.205 -26.935 17.345 -26.765 ;
      RECT 17.205 -25.439 17.295 -24.432 ;
      RECT 17.205 -24.915 17.345 -24.745 ;
      RECT 17.205 -24.018 17.295 -23.011 ;
      RECT 17.205 -23.705 17.345 -23.535 ;
      RECT 17.205 -22.209 17.295 -21.202 ;
      RECT 17.205 -21.685 17.345 -21.515 ;
      RECT 17.205 -20.788 17.295 -19.781 ;
      RECT 17.205 -20.475 17.345 -20.305 ;
      RECT 17.205 -18.979 17.295 -17.972 ;
      RECT 17.205 -18.455 17.345 -18.285 ;
      RECT 17.205 -17.558 17.295 -16.551 ;
      RECT 17.205 -17.245 17.345 -17.075 ;
      RECT 17.205 -15.749 17.295 -14.742 ;
      RECT 17.205 -15.225 17.345 -15.055 ;
      RECT 17.205 -14.328 17.295 -13.321 ;
      RECT 17.205 -14.015 17.345 -13.845 ;
      RECT 17.205 -12.519 17.295 -11.512 ;
      RECT 17.205 -11.995 17.345 -11.825 ;
      RECT 17.205 -11.098 17.295 -10.091 ;
      RECT 17.205 -10.785 17.345 -10.615 ;
      RECT 17.205 -9.289 17.295 -8.282 ;
      RECT 17.205 -8.765 17.345 -8.595 ;
      RECT 17.205 -7.868 17.295 -6.861 ;
      RECT 17.205 -7.555 17.345 -7.385 ;
      RECT 17.205 -6.059 17.295 -5.052 ;
      RECT 17.205 -5.535 17.345 -5.365 ;
      RECT 17.205 -4.638 17.295 -3.631 ;
      RECT 17.205 -4.325 17.345 -4.155 ;
      RECT 17.205 -2.829 17.295 -1.822 ;
      RECT 17.205 -2.305 17.345 -2.135 ;
      RECT 17.205 -1.408 17.295 -0.401 ;
      RECT 17.205 -1.095 17.345 -0.925 ;
      RECT 17.205 0.401 17.295 1.408 ;
      RECT 17.205 0.925 17.345 1.095 ;
      RECT 15.355 -60.005 16.835 -59.905 ;
      RECT 15.355 -60.375 15.455 -59.905 ;
      RECT 15.16 -62.715 16.735 -62.595 ;
      RECT 16.635 -63.215 16.735 -62.595 ;
      RECT 16.04 -63.215 16.14 -62.595 ;
      RECT 15.16 -63.17 15.26 -62.595 ;
      RECT 16.405 -49.858 16.495 -48.85 ;
      RECT 16.355 -49.255 16.495 -49.085 ;
      RECT 16.405 -48.05 16.495 -47.042 ;
      RECT 16.355 -47.815 16.495 -47.645 ;
      RECT 16.405 -46.628 16.495 -45.62 ;
      RECT 16.355 -46.025 16.495 -45.855 ;
      RECT 16.405 -44.82 16.495 -43.812 ;
      RECT 16.355 -44.585 16.495 -44.415 ;
      RECT 16.405 -43.398 16.495 -42.39 ;
      RECT 16.355 -42.795 16.495 -42.625 ;
      RECT 16.405 -41.59 16.495 -40.582 ;
      RECT 16.355 -41.355 16.495 -41.185 ;
      RECT 16.405 -40.168 16.495 -39.16 ;
      RECT 16.355 -39.565 16.495 -39.395 ;
      RECT 16.405 -38.36 16.495 -37.352 ;
      RECT 16.355 -38.125 16.495 -37.955 ;
      RECT 16.405 -36.938 16.495 -35.93 ;
      RECT 16.355 -36.335 16.495 -36.165 ;
      RECT 16.405 -35.13 16.495 -34.122 ;
      RECT 16.355 -34.895 16.495 -34.725 ;
      RECT 16.405 -33.708 16.495 -32.7 ;
      RECT 16.355 -33.105 16.495 -32.935 ;
      RECT 16.405 -31.9 16.495 -30.892 ;
      RECT 16.355 -31.665 16.495 -31.495 ;
      RECT 16.405 -30.478 16.495 -29.47 ;
      RECT 16.355 -29.875 16.495 -29.705 ;
      RECT 16.405 -28.67 16.495 -27.662 ;
      RECT 16.355 -28.435 16.495 -28.265 ;
      RECT 16.405 -27.248 16.495 -26.24 ;
      RECT 16.355 -26.645 16.495 -26.475 ;
      RECT 16.405 -25.44 16.495 -24.432 ;
      RECT 16.355 -25.205 16.495 -25.035 ;
      RECT 16.405 -24.018 16.495 -23.01 ;
      RECT 16.355 -23.415 16.495 -23.245 ;
      RECT 16.405 -22.21 16.495 -21.202 ;
      RECT 16.355 -21.975 16.495 -21.805 ;
      RECT 16.405 -20.788 16.495 -19.78 ;
      RECT 16.355 -20.185 16.495 -20.015 ;
      RECT 16.405 -18.98 16.495 -17.972 ;
      RECT 16.355 -18.745 16.495 -18.575 ;
      RECT 16.405 -17.558 16.495 -16.55 ;
      RECT 16.355 -16.955 16.495 -16.785 ;
      RECT 16.405 -15.75 16.495 -14.742 ;
      RECT 16.355 -15.515 16.495 -15.345 ;
      RECT 16.405 -14.328 16.495 -13.32 ;
      RECT 16.355 -13.725 16.495 -13.555 ;
      RECT 16.405 -12.52 16.495 -11.512 ;
      RECT 16.355 -12.285 16.495 -12.115 ;
      RECT 16.405 -11.098 16.495 -10.09 ;
      RECT 16.355 -10.495 16.495 -10.325 ;
      RECT 16.405 -9.29 16.495 -8.282 ;
      RECT 16.355 -9.055 16.495 -8.885 ;
      RECT 16.405 -7.868 16.495 -6.86 ;
      RECT 16.355 -7.265 16.495 -7.095 ;
      RECT 16.405 -6.06 16.495 -5.052 ;
      RECT 16.355 -5.825 16.495 -5.655 ;
      RECT 16.405 -4.638 16.495 -3.63 ;
      RECT 16.355 -4.035 16.495 -3.865 ;
      RECT 16.405 -2.83 16.495 -1.822 ;
      RECT 16.355 -2.595 16.495 -2.425 ;
      RECT 16.405 -1.408 16.495 -0.4 ;
      RECT 16.355 -0.805 16.495 -0.635 ;
      RECT 16.405 0.4 16.495 1.408 ;
      RECT 16.355 0.635 16.495 0.805 ;
      RECT 16.28 -63.005 16.455 -62.835 ;
      RECT 16.355 -63.215 16.455 -62.835 ;
      RECT 15.395 -61.875 15.495 -61.41 ;
      RECT 15.76 -61.875 15.86 -61.42 ;
      RECT 15.395 -61.875 16.24 -61.705 ;
      RECT 16.005 -49.858 16.095 -48.851 ;
      RECT 16.005 -49.545 16.145 -49.375 ;
      RECT 16.005 -48.049 16.095 -47.042 ;
      RECT 16.005 -47.525 16.145 -47.355 ;
      RECT 16.005 -46.628 16.095 -45.621 ;
      RECT 16.005 -46.315 16.145 -46.145 ;
      RECT 16.005 -44.819 16.095 -43.812 ;
      RECT 16.005 -44.295 16.145 -44.125 ;
      RECT 16.005 -43.398 16.095 -42.391 ;
      RECT 16.005 -43.085 16.145 -42.915 ;
      RECT 16.005 -41.589 16.095 -40.582 ;
      RECT 16.005 -41.065 16.145 -40.895 ;
      RECT 16.005 -40.168 16.095 -39.161 ;
      RECT 16.005 -39.855 16.145 -39.685 ;
      RECT 16.005 -38.359 16.095 -37.352 ;
      RECT 16.005 -37.835 16.145 -37.665 ;
      RECT 16.005 -36.938 16.095 -35.931 ;
      RECT 16.005 -36.625 16.145 -36.455 ;
      RECT 16.005 -35.129 16.095 -34.122 ;
      RECT 16.005 -34.605 16.145 -34.435 ;
      RECT 16.005 -33.708 16.095 -32.701 ;
      RECT 16.005 -33.395 16.145 -33.225 ;
      RECT 16.005 -31.899 16.095 -30.892 ;
      RECT 16.005 -31.375 16.145 -31.205 ;
      RECT 16.005 -30.478 16.095 -29.471 ;
      RECT 16.005 -30.165 16.145 -29.995 ;
      RECT 16.005 -28.669 16.095 -27.662 ;
      RECT 16.005 -28.145 16.145 -27.975 ;
      RECT 16.005 -27.248 16.095 -26.241 ;
      RECT 16.005 -26.935 16.145 -26.765 ;
      RECT 16.005 -25.439 16.095 -24.432 ;
      RECT 16.005 -24.915 16.145 -24.745 ;
      RECT 16.005 -24.018 16.095 -23.011 ;
      RECT 16.005 -23.705 16.145 -23.535 ;
      RECT 16.005 -22.209 16.095 -21.202 ;
      RECT 16.005 -21.685 16.145 -21.515 ;
      RECT 16.005 -20.788 16.095 -19.781 ;
      RECT 16.005 -20.475 16.145 -20.305 ;
      RECT 16.005 -18.979 16.095 -17.972 ;
      RECT 16.005 -18.455 16.145 -18.285 ;
      RECT 16.005 -17.558 16.095 -16.551 ;
      RECT 16.005 -17.245 16.145 -17.075 ;
      RECT 16.005 -15.749 16.095 -14.742 ;
      RECT 16.005 -15.225 16.145 -15.055 ;
      RECT 16.005 -14.328 16.095 -13.321 ;
      RECT 16.005 -14.015 16.145 -13.845 ;
      RECT 16.005 -12.519 16.095 -11.512 ;
      RECT 16.005 -11.995 16.145 -11.825 ;
      RECT 16.005 -11.098 16.095 -10.091 ;
      RECT 16.005 -10.785 16.145 -10.615 ;
      RECT 16.005 -9.289 16.095 -8.282 ;
      RECT 16.005 -8.765 16.145 -8.595 ;
      RECT 16.005 -7.868 16.095 -6.861 ;
      RECT 16.005 -7.555 16.145 -7.385 ;
      RECT 16.005 -6.059 16.095 -5.052 ;
      RECT 16.005 -5.535 16.145 -5.365 ;
      RECT 16.005 -4.638 16.095 -3.631 ;
      RECT 16.005 -4.325 16.145 -4.155 ;
      RECT 16.005 -2.829 16.095 -1.822 ;
      RECT 16.005 -2.305 16.145 -2.135 ;
      RECT 16.005 -1.408 16.095 -0.401 ;
      RECT 16.005 -1.095 16.145 -0.925 ;
      RECT 16.005 0.401 16.095 1.408 ;
      RECT 16.005 0.925 16.145 1.095 ;
      RECT 15.69 -63.005 15.86 -62.835 ;
      RECT 15.76 -63.215 15.86 -62.835 ;
      RECT 15.205 -49.858 15.295 -48.85 ;
      RECT 15.155 -49.255 15.295 -49.085 ;
      RECT 15.205 -48.05 15.295 -47.042 ;
      RECT 15.155 -47.815 15.295 -47.645 ;
      RECT 15.205 -46.628 15.295 -45.62 ;
      RECT 15.155 -46.025 15.295 -45.855 ;
      RECT 15.205 -44.82 15.295 -43.812 ;
      RECT 15.155 -44.585 15.295 -44.415 ;
      RECT 15.205 -43.398 15.295 -42.39 ;
      RECT 15.155 -42.795 15.295 -42.625 ;
      RECT 15.205 -41.59 15.295 -40.582 ;
      RECT 15.155 -41.355 15.295 -41.185 ;
      RECT 15.205 -40.168 15.295 -39.16 ;
      RECT 15.155 -39.565 15.295 -39.395 ;
      RECT 15.205 -38.36 15.295 -37.352 ;
      RECT 15.155 -38.125 15.295 -37.955 ;
      RECT 15.205 -36.938 15.295 -35.93 ;
      RECT 15.155 -36.335 15.295 -36.165 ;
      RECT 15.205 -35.13 15.295 -34.122 ;
      RECT 15.155 -34.895 15.295 -34.725 ;
      RECT 15.205 -33.708 15.295 -32.7 ;
      RECT 15.155 -33.105 15.295 -32.935 ;
      RECT 15.205 -31.9 15.295 -30.892 ;
      RECT 15.155 -31.665 15.295 -31.495 ;
      RECT 15.205 -30.478 15.295 -29.47 ;
      RECT 15.155 -29.875 15.295 -29.705 ;
      RECT 15.205 -28.67 15.295 -27.662 ;
      RECT 15.155 -28.435 15.295 -28.265 ;
      RECT 15.205 -27.248 15.295 -26.24 ;
      RECT 15.155 -26.645 15.295 -26.475 ;
      RECT 15.205 -25.44 15.295 -24.432 ;
      RECT 15.155 -25.205 15.295 -25.035 ;
      RECT 15.205 -24.018 15.295 -23.01 ;
      RECT 15.155 -23.415 15.295 -23.245 ;
      RECT 15.205 -22.21 15.295 -21.202 ;
      RECT 15.155 -21.975 15.295 -21.805 ;
      RECT 15.205 -20.788 15.295 -19.78 ;
      RECT 15.155 -20.185 15.295 -20.015 ;
      RECT 15.205 -18.98 15.295 -17.972 ;
      RECT 15.155 -18.745 15.295 -18.575 ;
      RECT 15.205 -17.558 15.295 -16.55 ;
      RECT 15.155 -16.955 15.295 -16.785 ;
      RECT 15.205 -15.75 15.295 -14.742 ;
      RECT 15.155 -15.515 15.295 -15.345 ;
      RECT 15.205 -14.328 15.295 -13.32 ;
      RECT 15.155 -13.725 15.295 -13.555 ;
      RECT 15.205 -12.52 15.295 -11.512 ;
      RECT 15.155 -12.285 15.295 -12.115 ;
      RECT 15.205 -11.098 15.295 -10.09 ;
      RECT 15.155 -10.495 15.295 -10.325 ;
      RECT 15.205 -9.29 15.295 -8.282 ;
      RECT 15.155 -9.055 15.295 -8.885 ;
      RECT 15.205 -7.868 15.295 -6.86 ;
      RECT 15.155 -7.265 15.295 -7.095 ;
      RECT 15.205 -6.06 15.295 -5.052 ;
      RECT 15.155 -5.825 15.295 -5.655 ;
      RECT 15.205 -4.638 15.295 -3.63 ;
      RECT 15.155 -4.035 15.295 -3.865 ;
      RECT 15.205 -2.83 15.295 -1.822 ;
      RECT 15.155 -2.595 15.295 -2.425 ;
      RECT 15.205 -1.408 15.295 -0.4 ;
      RECT 15.155 -0.805 15.295 -0.635 ;
      RECT 15.205 0.4 15.295 1.408 ;
      RECT 15.155 0.635 15.295 0.805 ;
      RECT 14.805 -49.858 14.895 -48.851 ;
      RECT 14.805 -49.545 14.945 -49.375 ;
      RECT 14.805 -48.049 14.895 -47.042 ;
      RECT 14.805 -47.525 14.945 -47.355 ;
      RECT 14.805 -46.628 14.895 -45.621 ;
      RECT 14.805 -46.315 14.945 -46.145 ;
      RECT 14.805 -44.819 14.895 -43.812 ;
      RECT 14.805 -44.295 14.945 -44.125 ;
      RECT 14.805 -43.398 14.895 -42.391 ;
      RECT 14.805 -43.085 14.945 -42.915 ;
      RECT 14.805 -41.589 14.895 -40.582 ;
      RECT 14.805 -41.065 14.945 -40.895 ;
      RECT 14.805 -40.168 14.895 -39.161 ;
      RECT 14.805 -39.855 14.945 -39.685 ;
      RECT 14.805 -38.359 14.895 -37.352 ;
      RECT 14.805 -37.835 14.945 -37.665 ;
      RECT 14.805 -36.938 14.895 -35.931 ;
      RECT 14.805 -36.625 14.945 -36.455 ;
      RECT 14.805 -35.129 14.895 -34.122 ;
      RECT 14.805 -34.605 14.945 -34.435 ;
      RECT 14.805 -33.708 14.895 -32.701 ;
      RECT 14.805 -33.395 14.945 -33.225 ;
      RECT 14.805 -31.899 14.895 -30.892 ;
      RECT 14.805 -31.375 14.945 -31.205 ;
      RECT 14.805 -30.478 14.895 -29.471 ;
      RECT 14.805 -30.165 14.945 -29.995 ;
      RECT 14.805 -28.669 14.895 -27.662 ;
      RECT 14.805 -28.145 14.945 -27.975 ;
      RECT 14.805 -27.248 14.895 -26.241 ;
      RECT 14.805 -26.935 14.945 -26.765 ;
      RECT 14.805 -25.439 14.895 -24.432 ;
      RECT 14.805 -24.915 14.945 -24.745 ;
      RECT 14.805 -24.018 14.895 -23.011 ;
      RECT 14.805 -23.705 14.945 -23.535 ;
      RECT 14.805 -22.209 14.895 -21.202 ;
      RECT 14.805 -21.685 14.945 -21.515 ;
      RECT 14.805 -20.788 14.895 -19.781 ;
      RECT 14.805 -20.475 14.945 -20.305 ;
      RECT 14.805 -18.979 14.895 -17.972 ;
      RECT 14.805 -18.455 14.945 -18.285 ;
      RECT 14.805 -17.558 14.895 -16.551 ;
      RECT 14.805 -17.245 14.945 -17.075 ;
      RECT 14.805 -15.749 14.895 -14.742 ;
      RECT 14.805 -15.225 14.945 -15.055 ;
      RECT 14.805 -14.328 14.895 -13.321 ;
      RECT 14.805 -14.015 14.945 -13.845 ;
      RECT 14.805 -12.519 14.895 -11.512 ;
      RECT 14.805 -11.995 14.945 -11.825 ;
      RECT 14.805 -11.098 14.895 -10.091 ;
      RECT 14.805 -10.785 14.945 -10.615 ;
      RECT 14.805 -9.289 14.895 -8.282 ;
      RECT 14.805 -8.765 14.945 -8.595 ;
      RECT 14.805 -7.868 14.895 -6.861 ;
      RECT 14.805 -7.555 14.945 -7.385 ;
      RECT 14.805 -6.059 14.895 -5.052 ;
      RECT 14.805 -5.535 14.945 -5.365 ;
      RECT 14.805 -4.638 14.895 -3.631 ;
      RECT 14.805 -4.325 14.945 -4.155 ;
      RECT 14.805 -2.829 14.895 -1.822 ;
      RECT 14.805 -2.305 14.945 -2.135 ;
      RECT 14.805 -1.408 14.895 -0.401 ;
      RECT 14.805 -1.095 14.945 -0.925 ;
      RECT 14.805 0.401 14.895 1.408 ;
      RECT 14.805 0.925 14.945 1.095 ;
      RECT 10.635 -57.255 14.415 -57.135 ;
      RECT 11.955 -57.795 12.055 -57.135 ;
      RECT 11.395 -57.795 11.495 -57.135 ;
      RECT 10.835 -57.795 10.935 -57.135 ;
      RECT 14.005 -49.858 14.095 -48.85 ;
      RECT 13.955 -49.255 14.095 -49.085 ;
      RECT 14.005 -48.05 14.095 -47.042 ;
      RECT 13.955 -47.815 14.095 -47.645 ;
      RECT 14.005 -46.628 14.095 -45.62 ;
      RECT 13.955 -46.025 14.095 -45.855 ;
      RECT 14.005 -44.82 14.095 -43.812 ;
      RECT 13.955 -44.585 14.095 -44.415 ;
      RECT 14.005 -43.398 14.095 -42.39 ;
      RECT 13.955 -42.795 14.095 -42.625 ;
      RECT 14.005 -41.59 14.095 -40.582 ;
      RECT 13.955 -41.355 14.095 -41.185 ;
      RECT 14.005 -40.168 14.095 -39.16 ;
      RECT 13.955 -39.565 14.095 -39.395 ;
      RECT 14.005 -38.36 14.095 -37.352 ;
      RECT 13.955 -38.125 14.095 -37.955 ;
      RECT 14.005 -36.938 14.095 -35.93 ;
      RECT 13.955 -36.335 14.095 -36.165 ;
      RECT 14.005 -35.13 14.095 -34.122 ;
      RECT 13.955 -34.895 14.095 -34.725 ;
      RECT 14.005 -33.708 14.095 -32.7 ;
      RECT 13.955 -33.105 14.095 -32.935 ;
      RECT 14.005 -31.9 14.095 -30.892 ;
      RECT 13.955 -31.665 14.095 -31.495 ;
      RECT 14.005 -30.478 14.095 -29.47 ;
      RECT 13.955 -29.875 14.095 -29.705 ;
      RECT 14.005 -28.67 14.095 -27.662 ;
      RECT 13.955 -28.435 14.095 -28.265 ;
      RECT 14.005 -27.248 14.095 -26.24 ;
      RECT 13.955 -26.645 14.095 -26.475 ;
      RECT 14.005 -25.44 14.095 -24.432 ;
      RECT 13.955 -25.205 14.095 -25.035 ;
      RECT 14.005 -24.018 14.095 -23.01 ;
      RECT 13.955 -23.415 14.095 -23.245 ;
      RECT 14.005 -22.21 14.095 -21.202 ;
      RECT 13.955 -21.975 14.095 -21.805 ;
      RECT 14.005 -20.788 14.095 -19.78 ;
      RECT 13.955 -20.185 14.095 -20.015 ;
      RECT 14.005 -18.98 14.095 -17.972 ;
      RECT 13.955 -18.745 14.095 -18.575 ;
      RECT 14.005 -17.558 14.095 -16.55 ;
      RECT 13.955 -16.955 14.095 -16.785 ;
      RECT 14.005 -15.75 14.095 -14.742 ;
      RECT 13.955 -15.515 14.095 -15.345 ;
      RECT 14.005 -14.328 14.095 -13.32 ;
      RECT 13.955 -13.725 14.095 -13.555 ;
      RECT 14.005 -12.52 14.095 -11.512 ;
      RECT 13.955 -12.285 14.095 -12.115 ;
      RECT 14.005 -11.098 14.095 -10.09 ;
      RECT 13.955 -10.495 14.095 -10.325 ;
      RECT 14.005 -9.29 14.095 -8.282 ;
      RECT 13.955 -9.055 14.095 -8.885 ;
      RECT 14.005 -7.868 14.095 -6.86 ;
      RECT 13.955 -7.265 14.095 -7.095 ;
      RECT 14.005 -6.06 14.095 -5.052 ;
      RECT 13.955 -5.825 14.095 -5.655 ;
      RECT 14.005 -4.638 14.095 -3.63 ;
      RECT 13.955 -4.035 14.095 -3.865 ;
      RECT 14.005 -2.83 14.095 -1.822 ;
      RECT 13.955 -2.595 14.095 -2.425 ;
      RECT 14.005 -1.408 14.095 -0.4 ;
      RECT 13.955 -0.805 14.095 -0.635 ;
      RECT 14.005 0.4 14.095 1.408 ;
      RECT 13.955 0.635 14.095 0.805 ;
      RECT 12.575 -60.005 14.055 -59.905 ;
      RECT 12.575 -60.515 12.675 -59.905 ;
      RECT 12.795 -57.47 14.055 -57.37 ;
      RECT 13.955 -57.795 14.055 -57.37 ;
      RECT 13.395 -57.795 13.495 -57.37 ;
      RECT 12.835 -57.795 12.935 -57.37 ;
      RECT 13.605 -49.858 13.695 -48.851 ;
      RECT 13.605 -49.545 13.745 -49.375 ;
      RECT 13.605 -48.049 13.695 -47.042 ;
      RECT 13.605 -47.525 13.745 -47.355 ;
      RECT 13.605 -46.628 13.695 -45.621 ;
      RECT 13.605 -46.315 13.745 -46.145 ;
      RECT 13.605 -44.819 13.695 -43.812 ;
      RECT 13.605 -44.295 13.745 -44.125 ;
      RECT 13.605 -43.398 13.695 -42.391 ;
      RECT 13.605 -43.085 13.745 -42.915 ;
      RECT 13.605 -41.589 13.695 -40.582 ;
      RECT 13.605 -41.065 13.745 -40.895 ;
      RECT 13.605 -40.168 13.695 -39.161 ;
      RECT 13.605 -39.855 13.745 -39.685 ;
      RECT 13.605 -38.359 13.695 -37.352 ;
      RECT 13.605 -37.835 13.745 -37.665 ;
      RECT 13.605 -36.938 13.695 -35.931 ;
      RECT 13.605 -36.625 13.745 -36.455 ;
      RECT 13.605 -35.129 13.695 -34.122 ;
      RECT 13.605 -34.605 13.745 -34.435 ;
      RECT 13.605 -33.708 13.695 -32.701 ;
      RECT 13.605 -33.395 13.745 -33.225 ;
      RECT 13.605 -31.899 13.695 -30.892 ;
      RECT 13.605 -31.375 13.745 -31.205 ;
      RECT 13.605 -30.478 13.695 -29.471 ;
      RECT 13.605 -30.165 13.745 -29.995 ;
      RECT 13.605 -28.669 13.695 -27.662 ;
      RECT 13.605 -28.145 13.745 -27.975 ;
      RECT 13.605 -27.248 13.695 -26.241 ;
      RECT 13.605 -26.935 13.745 -26.765 ;
      RECT 13.605 -25.439 13.695 -24.432 ;
      RECT 13.605 -24.915 13.745 -24.745 ;
      RECT 13.605 -24.018 13.695 -23.011 ;
      RECT 13.605 -23.705 13.745 -23.535 ;
      RECT 13.605 -22.209 13.695 -21.202 ;
      RECT 13.605 -21.685 13.745 -21.515 ;
      RECT 13.605 -20.788 13.695 -19.781 ;
      RECT 13.605 -20.475 13.745 -20.305 ;
      RECT 13.605 -18.979 13.695 -17.972 ;
      RECT 13.605 -18.455 13.745 -18.285 ;
      RECT 13.605 -17.558 13.695 -16.551 ;
      RECT 13.605 -17.245 13.745 -17.075 ;
      RECT 13.605 -15.749 13.695 -14.742 ;
      RECT 13.605 -15.225 13.745 -15.055 ;
      RECT 13.605 -14.328 13.695 -13.321 ;
      RECT 13.605 -14.015 13.745 -13.845 ;
      RECT 13.605 -12.519 13.695 -11.512 ;
      RECT 13.605 -11.995 13.745 -11.825 ;
      RECT 13.605 -11.098 13.695 -10.091 ;
      RECT 13.605 -10.785 13.745 -10.615 ;
      RECT 13.605 -9.289 13.695 -8.282 ;
      RECT 13.605 -8.765 13.745 -8.595 ;
      RECT 13.605 -7.868 13.695 -6.861 ;
      RECT 13.605 -7.555 13.745 -7.385 ;
      RECT 13.605 -6.059 13.695 -5.052 ;
      RECT 13.605 -5.535 13.745 -5.365 ;
      RECT 13.605 -4.638 13.695 -3.631 ;
      RECT 13.605 -4.325 13.745 -4.155 ;
      RECT 13.605 -2.829 13.695 -1.822 ;
      RECT 13.605 -2.305 13.745 -2.135 ;
      RECT 13.605 -1.408 13.695 -0.401 ;
      RECT 13.605 -1.095 13.745 -0.925 ;
      RECT 13.605 0.401 13.695 1.408 ;
      RECT 13.605 0.925 13.745 1.095 ;
      RECT 12.935 -59.815 13.105 -59.705 ;
      RECT 9.785 -59.815 13.105 -59.715 ;
      RECT 12.805 -49.858 12.895 -48.85 ;
      RECT 12.755 -49.255 12.895 -49.085 ;
      RECT 12.805 -48.05 12.895 -47.042 ;
      RECT 12.755 -47.815 12.895 -47.645 ;
      RECT 12.805 -46.628 12.895 -45.62 ;
      RECT 12.755 -46.025 12.895 -45.855 ;
      RECT 12.805 -44.82 12.895 -43.812 ;
      RECT 12.755 -44.585 12.895 -44.415 ;
      RECT 12.805 -43.398 12.895 -42.39 ;
      RECT 12.755 -42.795 12.895 -42.625 ;
      RECT 12.805 -41.59 12.895 -40.582 ;
      RECT 12.755 -41.355 12.895 -41.185 ;
      RECT 12.805 -40.168 12.895 -39.16 ;
      RECT 12.755 -39.565 12.895 -39.395 ;
      RECT 12.805 -38.36 12.895 -37.352 ;
      RECT 12.755 -38.125 12.895 -37.955 ;
      RECT 12.805 -36.938 12.895 -35.93 ;
      RECT 12.755 -36.335 12.895 -36.165 ;
      RECT 12.805 -35.13 12.895 -34.122 ;
      RECT 12.755 -34.895 12.895 -34.725 ;
      RECT 12.805 -33.708 12.895 -32.7 ;
      RECT 12.755 -33.105 12.895 -32.935 ;
      RECT 12.805 -31.9 12.895 -30.892 ;
      RECT 12.755 -31.665 12.895 -31.495 ;
      RECT 12.805 -30.478 12.895 -29.47 ;
      RECT 12.755 -29.875 12.895 -29.705 ;
      RECT 12.805 -28.67 12.895 -27.662 ;
      RECT 12.755 -28.435 12.895 -28.265 ;
      RECT 12.805 -27.248 12.895 -26.24 ;
      RECT 12.755 -26.645 12.895 -26.475 ;
      RECT 12.805 -25.44 12.895 -24.432 ;
      RECT 12.755 -25.205 12.895 -25.035 ;
      RECT 12.805 -24.018 12.895 -23.01 ;
      RECT 12.755 -23.415 12.895 -23.245 ;
      RECT 12.805 -22.21 12.895 -21.202 ;
      RECT 12.755 -21.975 12.895 -21.805 ;
      RECT 12.805 -20.788 12.895 -19.78 ;
      RECT 12.755 -20.185 12.895 -20.015 ;
      RECT 12.805 -18.98 12.895 -17.972 ;
      RECT 12.755 -18.745 12.895 -18.575 ;
      RECT 12.805 -17.558 12.895 -16.55 ;
      RECT 12.755 -16.955 12.895 -16.785 ;
      RECT 12.805 -15.75 12.895 -14.742 ;
      RECT 12.755 -15.515 12.895 -15.345 ;
      RECT 12.805 -14.328 12.895 -13.32 ;
      RECT 12.755 -13.725 12.895 -13.555 ;
      RECT 12.805 -12.52 12.895 -11.512 ;
      RECT 12.755 -12.285 12.895 -12.115 ;
      RECT 12.805 -11.098 12.895 -10.09 ;
      RECT 12.755 -10.495 12.895 -10.325 ;
      RECT 12.805 -9.29 12.895 -8.282 ;
      RECT 12.755 -9.055 12.895 -8.885 ;
      RECT 12.805 -7.868 12.895 -6.86 ;
      RECT 12.755 -7.265 12.895 -7.095 ;
      RECT 12.805 -6.06 12.895 -5.052 ;
      RECT 12.755 -5.825 12.895 -5.655 ;
      RECT 12.805 -4.638 12.895 -3.63 ;
      RECT 12.755 -4.035 12.895 -3.865 ;
      RECT 12.805 -2.83 12.895 -1.822 ;
      RECT 12.755 -2.595 12.895 -2.425 ;
      RECT 12.805 -1.408 12.895 -0.4 ;
      RECT 12.755 -0.805 12.895 -0.635 ;
      RECT 12.805 0.4 12.895 1.408 ;
      RECT 12.755 0.635 12.895 0.805 ;
      RECT 12.405 -49.858 12.495 -48.851 ;
      RECT 12.405 -49.545 12.545 -49.375 ;
      RECT 12.405 -48.049 12.495 -47.042 ;
      RECT 12.405 -47.525 12.545 -47.355 ;
      RECT 12.405 -46.628 12.495 -45.621 ;
      RECT 12.405 -46.315 12.545 -46.145 ;
      RECT 12.405 -44.819 12.495 -43.812 ;
      RECT 12.405 -44.295 12.545 -44.125 ;
      RECT 12.405 -43.398 12.495 -42.391 ;
      RECT 12.405 -43.085 12.545 -42.915 ;
      RECT 12.405 -41.589 12.495 -40.582 ;
      RECT 12.405 -41.065 12.545 -40.895 ;
      RECT 12.405 -40.168 12.495 -39.161 ;
      RECT 12.405 -39.855 12.545 -39.685 ;
      RECT 12.405 -38.359 12.495 -37.352 ;
      RECT 12.405 -37.835 12.545 -37.665 ;
      RECT 12.405 -36.938 12.495 -35.931 ;
      RECT 12.405 -36.625 12.545 -36.455 ;
      RECT 12.405 -35.129 12.495 -34.122 ;
      RECT 12.405 -34.605 12.545 -34.435 ;
      RECT 12.405 -33.708 12.495 -32.701 ;
      RECT 12.405 -33.395 12.545 -33.225 ;
      RECT 12.405 -31.899 12.495 -30.892 ;
      RECT 12.405 -31.375 12.545 -31.205 ;
      RECT 12.405 -30.478 12.495 -29.471 ;
      RECT 12.405 -30.165 12.545 -29.995 ;
      RECT 12.405 -28.669 12.495 -27.662 ;
      RECT 12.405 -28.145 12.545 -27.975 ;
      RECT 12.405 -27.248 12.495 -26.241 ;
      RECT 12.405 -26.935 12.545 -26.765 ;
      RECT 12.405 -25.439 12.495 -24.432 ;
      RECT 12.405 -24.915 12.545 -24.745 ;
      RECT 12.405 -24.018 12.495 -23.011 ;
      RECT 12.405 -23.705 12.545 -23.535 ;
      RECT 12.405 -22.209 12.495 -21.202 ;
      RECT 12.405 -21.685 12.545 -21.515 ;
      RECT 12.405 -20.788 12.495 -19.781 ;
      RECT 12.405 -20.475 12.545 -20.305 ;
      RECT 12.405 -18.979 12.495 -17.972 ;
      RECT 12.405 -18.455 12.545 -18.285 ;
      RECT 12.405 -17.558 12.495 -16.551 ;
      RECT 12.405 -17.245 12.545 -17.075 ;
      RECT 12.405 -15.749 12.495 -14.742 ;
      RECT 12.405 -15.225 12.545 -15.055 ;
      RECT 12.405 -14.328 12.495 -13.321 ;
      RECT 12.405 -14.015 12.545 -13.845 ;
      RECT 12.405 -12.519 12.495 -11.512 ;
      RECT 12.405 -11.995 12.545 -11.825 ;
      RECT 12.405 -11.098 12.495 -10.091 ;
      RECT 12.405 -10.785 12.545 -10.615 ;
      RECT 12.405 -9.289 12.495 -8.282 ;
      RECT 12.405 -8.765 12.545 -8.595 ;
      RECT 12.405 -7.868 12.495 -6.861 ;
      RECT 12.405 -7.555 12.545 -7.385 ;
      RECT 12.405 -6.059 12.495 -5.052 ;
      RECT 12.405 -5.535 12.545 -5.365 ;
      RECT 12.405 -4.638 12.495 -3.631 ;
      RECT 12.405 -4.325 12.545 -4.155 ;
      RECT 12.405 -2.829 12.495 -1.822 ;
      RECT 12.405 -2.305 12.545 -2.135 ;
      RECT 12.405 -1.408 12.495 -0.401 ;
      RECT 12.405 -1.095 12.545 -0.925 ;
      RECT 12.405 0.401 12.495 1.408 ;
      RECT 12.405 0.925 12.545 1.095 ;
      RECT 10.555 -60.005 12.035 -59.905 ;
      RECT 10.555 -60.375 10.655 -59.905 ;
      RECT 10.36 -62.715 11.935 -62.595 ;
      RECT 11.835 -63.215 11.935 -62.595 ;
      RECT 11.24 -63.215 11.34 -62.595 ;
      RECT 10.36 -63.17 10.46 -62.595 ;
      RECT 11.605 -49.858 11.695 -48.85 ;
      RECT 11.555 -49.255 11.695 -49.085 ;
      RECT 11.605 -48.05 11.695 -47.042 ;
      RECT 11.555 -47.815 11.695 -47.645 ;
      RECT 11.605 -46.628 11.695 -45.62 ;
      RECT 11.555 -46.025 11.695 -45.855 ;
      RECT 11.605 -44.82 11.695 -43.812 ;
      RECT 11.555 -44.585 11.695 -44.415 ;
      RECT 11.605 -43.398 11.695 -42.39 ;
      RECT 11.555 -42.795 11.695 -42.625 ;
      RECT 11.605 -41.59 11.695 -40.582 ;
      RECT 11.555 -41.355 11.695 -41.185 ;
      RECT 11.605 -40.168 11.695 -39.16 ;
      RECT 11.555 -39.565 11.695 -39.395 ;
      RECT 11.605 -38.36 11.695 -37.352 ;
      RECT 11.555 -38.125 11.695 -37.955 ;
      RECT 11.605 -36.938 11.695 -35.93 ;
      RECT 11.555 -36.335 11.695 -36.165 ;
      RECT 11.605 -35.13 11.695 -34.122 ;
      RECT 11.555 -34.895 11.695 -34.725 ;
      RECT 11.605 -33.708 11.695 -32.7 ;
      RECT 11.555 -33.105 11.695 -32.935 ;
      RECT 11.605 -31.9 11.695 -30.892 ;
      RECT 11.555 -31.665 11.695 -31.495 ;
      RECT 11.605 -30.478 11.695 -29.47 ;
      RECT 11.555 -29.875 11.695 -29.705 ;
      RECT 11.605 -28.67 11.695 -27.662 ;
      RECT 11.555 -28.435 11.695 -28.265 ;
      RECT 11.605 -27.248 11.695 -26.24 ;
      RECT 11.555 -26.645 11.695 -26.475 ;
      RECT 11.605 -25.44 11.695 -24.432 ;
      RECT 11.555 -25.205 11.695 -25.035 ;
      RECT 11.605 -24.018 11.695 -23.01 ;
      RECT 11.555 -23.415 11.695 -23.245 ;
      RECT 11.605 -22.21 11.695 -21.202 ;
      RECT 11.555 -21.975 11.695 -21.805 ;
      RECT 11.605 -20.788 11.695 -19.78 ;
      RECT 11.555 -20.185 11.695 -20.015 ;
      RECT 11.605 -18.98 11.695 -17.972 ;
      RECT 11.555 -18.745 11.695 -18.575 ;
      RECT 11.605 -17.558 11.695 -16.55 ;
      RECT 11.555 -16.955 11.695 -16.785 ;
      RECT 11.605 -15.75 11.695 -14.742 ;
      RECT 11.555 -15.515 11.695 -15.345 ;
      RECT 11.605 -14.328 11.695 -13.32 ;
      RECT 11.555 -13.725 11.695 -13.555 ;
      RECT 11.605 -12.52 11.695 -11.512 ;
      RECT 11.555 -12.285 11.695 -12.115 ;
      RECT 11.605 -11.098 11.695 -10.09 ;
      RECT 11.555 -10.495 11.695 -10.325 ;
      RECT 11.605 -9.29 11.695 -8.282 ;
      RECT 11.555 -9.055 11.695 -8.885 ;
      RECT 11.605 -7.868 11.695 -6.86 ;
      RECT 11.555 -7.265 11.695 -7.095 ;
      RECT 11.605 -6.06 11.695 -5.052 ;
      RECT 11.555 -5.825 11.695 -5.655 ;
      RECT 11.605 -4.638 11.695 -3.63 ;
      RECT 11.555 -4.035 11.695 -3.865 ;
      RECT 11.605 -2.83 11.695 -1.822 ;
      RECT 11.555 -2.595 11.695 -2.425 ;
      RECT 11.605 -1.408 11.695 -0.4 ;
      RECT 11.555 -0.805 11.695 -0.635 ;
      RECT 11.605 0.4 11.695 1.408 ;
      RECT 11.555 0.635 11.695 0.805 ;
      RECT 11.48 -63.005 11.655 -62.835 ;
      RECT 11.555 -63.215 11.655 -62.835 ;
      RECT 10.595 -61.875 10.695 -61.41 ;
      RECT 10.96 -61.875 11.06 -61.42 ;
      RECT 10.595 -61.875 11.44 -61.705 ;
      RECT 11.205 -49.858 11.295 -48.851 ;
      RECT 11.205 -49.545 11.345 -49.375 ;
      RECT 11.205 -48.049 11.295 -47.042 ;
      RECT 11.205 -47.525 11.345 -47.355 ;
      RECT 11.205 -46.628 11.295 -45.621 ;
      RECT 11.205 -46.315 11.345 -46.145 ;
      RECT 11.205 -44.819 11.295 -43.812 ;
      RECT 11.205 -44.295 11.345 -44.125 ;
      RECT 11.205 -43.398 11.295 -42.391 ;
      RECT 11.205 -43.085 11.345 -42.915 ;
      RECT 11.205 -41.589 11.295 -40.582 ;
      RECT 11.205 -41.065 11.345 -40.895 ;
      RECT 11.205 -40.168 11.295 -39.161 ;
      RECT 11.205 -39.855 11.345 -39.685 ;
      RECT 11.205 -38.359 11.295 -37.352 ;
      RECT 11.205 -37.835 11.345 -37.665 ;
      RECT 11.205 -36.938 11.295 -35.931 ;
      RECT 11.205 -36.625 11.345 -36.455 ;
      RECT 11.205 -35.129 11.295 -34.122 ;
      RECT 11.205 -34.605 11.345 -34.435 ;
      RECT 11.205 -33.708 11.295 -32.701 ;
      RECT 11.205 -33.395 11.345 -33.225 ;
      RECT 11.205 -31.899 11.295 -30.892 ;
      RECT 11.205 -31.375 11.345 -31.205 ;
      RECT 11.205 -30.478 11.295 -29.471 ;
      RECT 11.205 -30.165 11.345 -29.995 ;
      RECT 11.205 -28.669 11.295 -27.662 ;
      RECT 11.205 -28.145 11.345 -27.975 ;
      RECT 11.205 -27.248 11.295 -26.241 ;
      RECT 11.205 -26.935 11.345 -26.765 ;
      RECT 11.205 -25.439 11.295 -24.432 ;
      RECT 11.205 -24.915 11.345 -24.745 ;
      RECT 11.205 -24.018 11.295 -23.011 ;
      RECT 11.205 -23.705 11.345 -23.535 ;
      RECT 11.205 -22.209 11.295 -21.202 ;
      RECT 11.205 -21.685 11.345 -21.515 ;
      RECT 11.205 -20.788 11.295 -19.781 ;
      RECT 11.205 -20.475 11.345 -20.305 ;
      RECT 11.205 -18.979 11.295 -17.972 ;
      RECT 11.205 -18.455 11.345 -18.285 ;
      RECT 11.205 -17.558 11.295 -16.551 ;
      RECT 11.205 -17.245 11.345 -17.075 ;
      RECT 11.205 -15.749 11.295 -14.742 ;
      RECT 11.205 -15.225 11.345 -15.055 ;
      RECT 11.205 -14.328 11.295 -13.321 ;
      RECT 11.205 -14.015 11.345 -13.845 ;
      RECT 11.205 -12.519 11.295 -11.512 ;
      RECT 11.205 -11.995 11.345 -11.825 ;
      RECT 11.205 -11.098 11.295 -10.091 ;
      RECT 11.205 -10.785 11.345 -10.615 ;
      RECT 11.205 -9.289 11.295 -8.282 ;
      RECT 11.205 -8.765 11.345 -8.595 ;
      RECT 11.205 -7.868 11.295 -6.861 ;
      RECT 11.205 -7.555 11.345 -7.385 ;
      RECT 11.205 -6.059 11.295 -5.052 ;
      RECT 11.205 -5.535 11.345 -5.365 ;
      RECT 11.205 -4.638 11.295 -3.631 ;
      RECT 11.205 -4.325 11.345 -4.155 ;
      RECT 11.205 -2.829 11.295 -1.822 ;
      RECT 11.205 -2.305 11.345 -2.135 ;
      RECT 11.205 -1.408 11.295 -0.401 ;
      RECT 11.205 -1.095 11.345 -0.925 ;
      RECT 11.205 0.401 11.295 1.408 ;
      RECT 11.205 0.925 11.345 1.095 ;
      RECT 10.89 -63.005 11.06 -62.835 ;
      RECT 10.96 -63.215 11.06 -62.835 ;
      RECT 10.405 -49.858 10.495 -48.85 ;
      RECT 10.355 -49.255 10.495 -49.085 ;
      RECT 10.405 -48.05 10.495 -47.042 ;
      RECT 10.355 -47.815 10.495 -47.645 ;
      RECT 10.405 -46.628 10.495 -45.62 ;
      RECT 10.355 -46.025 10.495 -45.855 ;
      RECT 10.405 -44.82 10.495 -43.812 ;
      RECT 10.355 -44.585 10.495 -44.415 ;
      RECT 10.405 -43.398 10.495 -42.39 ;
      RECT 10.355 -42.795 10.495 -42.625 ;
      RECT 10.405 -41.59 10.495 -40.582 ;
      RECT 10.355 -41.355 10.495 -41.185 ;
      RECT 10.405 -40.168 10.495 -39.16 ;
      RECT 10.355 -39.565 10.495 -39.395 ;
      RECT 10.405 -38.36 10.495 -37.352 ;
      RECT 10.355 -38.125 10.495 -37.955 ;
      RECT 10.405 -36.938 10.495 -35.93 ;
      RECT 10.355 -36.335 10.495 -36.165 ;
      RECT 10.405 -35.13 10.495 -34.122 ;
      RECT 10.355 -34.895 10.495 -34.725 ;
      RECT 10.405 -33.708 10.495 -32.7 ;
      RECT 10.355 -33.105 10.495 -32.935 ;
      RECT 10.405 -31.9 10.495 -30.892 ;
      RECT 10.355 -31.665 10.495 -31.495 ;
      RECT 10.405 -30.478 10.495 -29.47 ;
      RECT 10.355 -29.875 10.495 -29.705 ;
      RECT 10.405 -28.67 10.495 -27.662 ;
      RECT 10.355 -28.435 10.495 -28.265 ;
      RECT 10.405 -27.248 10.495 -26.24 ;
      RECT 10.355 -26.645 10.495 -26.475 ;
      RECT 10.405 -25.44 10.495 -24.432 ;
      RECT 10.355 -25.205 10.495 -25.035 ;
      RECT 10.405 -24.018 10.495 -23.01 ;
      RECT 10.355 -23.415 10.495 -23.245 ;
      RECT 10.405 -22.21 10.495 -21.202 ;
      RECT 10.355 -21.975 10.495 -21.805 ;
      RECT 10.405 -20.788 10.495 -19.78 ;
      RECT 10.355 -20.185 10.495 -20.015 ;
      RECT 10.405 -18.98 10.495 -17.972 ;
      RECT 10.355 -18.745 10.495 -18.575 ;
      RECT 10.405 -17.558 10.495 -16.55 ;
      RECT 10.355 -16.955 10.495 -16.785 ;
      RECT 10.405 -15.75 10.495 -14.742 ;
      RECT 10.355 -15.515 10.495 -15.345 ;
      RECT 10.405 -14.328 10.495 -13.32 ;
      RECT 10.355 -13.725 10.495 -13.555 ;
      RECT 10.405 -12.52 10.495 -11.512 ;
      RECT 10.355 -12.285 10.495 -12.115 ;
      RECT 10.405 -11.098 10.495 -10.09 ;
      RECT 10.355 -10.495 10.495 -10.325 ;
      RECT 10.405 -9.29 10.495 -8.282 ;
      RECT 10.355 -9.055 10.495 -8.885 ;
      RECT 10.405 -7.868 10.495 -6.86 ;
      RECT 10.355 -7.265 10.495 -7.095 ;
      RECT 10.405 -6.06 10.495 -5.052 ;
      RECT 10.355 -5.825 10.495 -5.655 ;
      RECT 10.405 -4.638 10.495 -3.63 ;
      RECT 10.355 -4.035 10.495 -3.865 ;
      RECT 10.405 -2.83 10.495 -1.822 ;
      RECT 10.355 -2.595 10.495 -2.425 ;
      RECT 10.405 -1.408 10.495 -0.4 ;
      RECT 10.355 -0.805 10.495 -0.635 ;
      RECT 10.405 0.4 10.495 1.408 ;
      RECT 10.355 0.635 10.495 0.805 ;
      RECT 10.005 -49.858 10.095 -48.851 ;
      RECT 10.005 -49.545 10.145 -49.375 ;
      RECT 10.005 -48.049 10.095 -47.042 ;
      RECT 10.005 -47.525 10.145 -47.355 ;
      RECT 10.005 -46.628 10.095 -45.621 ;
      RECT 10.005 -46.315 10.145 -46.145 ;
      RECT 10.005 -44.819 10.095 -43.812 ;
      RECT 10.005 -44.295 10.145 -44.125 ;
      RECT 10.005 -43.398 10.095 -42.391 ;
      RECT 10.005 -43.085 10.145 -42.915 ;
      RECT 10.005 -41.589 10.095 -40.582 ;
      RECT 10.005 -41.065 10.145 -40.895 ;
      RECT 10.005 -40.168 10.095 -39.161 ;
      RECT 10.005 -39.855 10.145 -39.685 ;
      RECT 10.005 -38.359 10.095 -37.352 ;
      RECT 10.005 -37.835 10.145 -37.665 ;
      RECT 10.005 -36.938 10.095 -35.931 ;
      RECT 10.005 -36.625 10.145 -36.455 ;
      RECT 10.005 -35.129 10.095 -34.122 ;
      RECT 10.005 -34.605 10.145 -34.435 ;
      RECT 10.005 -33.708 10.095 -32.701 ;
      RECT 10.005 -33.395 10.145 -33.225 ;
      RECT 10.005 -31.899 10.095 -30.892 ;
      RECT 10.005 -31.375 10.145 -31.205 ;
      RECT 10.005 -30.478 10.095 -29.471 ;
      RECT 10.005 -30.165 10.145 -29.995 ;
      RECT 10.005 -28.669 10.095 -27.662 ;
      RECT 10.005 -28.145 10.145 -27.975 ;
      RECT 10.005 -27.248 10.095 -26.241 ;
      RECT 10.005 -26.935 10.145 -26.765 ;
      RECT 10.005 -25.439 10.095 -24.432 ;
      RECT 10.005 -24.915 10.145 -24.745 ;
      RECT 10.005 -24.018 10.095 -23.011 ;
      RECT 10.005 -23.705 10.145 -23.535 ;
      RECT 10.005 -22.209 10.095 -21.202 ;
      RECT 10.005 -21.685 10.145 -21.515 ;
      RECT 10.005 -20.788 10.095 -19.781 ;
      RECT 10.005 -20.475 10.145 -20.305 ;
      RECT 10.005 -18.979 10.095 -17.972 ;
      RECT 10.005 -18.455 10.145 -18.285 ;
      RECT 10.005 -17.558 10.095 -16.551 ;
      RECT 10.005 -17.245 10.145 -17.075 ;
      RECT 10.005 -15.749 10.095 -14.742 ;
      RECT 10.005 -15.225 10.145 -15.055 ;
      RECT 10.005 -14.328 10.095 -13.321 ;
      RECT 10.005 -14.015 10.145 -13.845 ;
      RECT 10.005 -12.519 10.095 -11.512 ;
      RECT 10.005 -11.995 10.145 -11.825 ;
      RECT 10.005 -11.098 10.095 -10.091 ;
      RECT 10.005 -10.785 10.145 -10.615 ;
      RECT 10.005 -9.289 10.095 -8.282 ;
      RECT 10.005 -8.765 10.145 -8.595 ;
      RECT 10.005 -7.868 10.095 -6.861 ;
      RECT 10.005 -7.555 10.145 -7.385 ;
      RECT 10.005 -6.059 10.095 -5.052 ;
      RECT 10.005 -5.535 10.145 -5.365 ;
      RECT 10.005 -4.638 10.095 -3.631 ;
      RECT 10.005 -4.325 10.145 -4.155 ;
      RECT 10.005 -2.829 10.095 -1.822 ;
      RECT 10.005 -2.305 10.145 -2.135 ;
      RECT 10.005 -1.408 10.095 -0.401 ;
      RECT 10.005 -1.095 10.145 -0.925 ;
      RECT 10.005 0.401 10.095 1.408 ;
      RECT 10.005 0.925 10.145 1.095 ;
      RECT 5.835 -57.255 9.615 -57.135 ;
      RECT 7.155 -57.795 7.255 -57.135 ;
      RECT 6.595 -57.795 6.695 -57.135 ;
      RECT 6.035 -57.795 6.135 -57.135 ;
      RECT 9.205 -49.858 9.295 -48.85 ;
      RECT 9.155 -49.255 9.295 -49.085 ;
      RECT 9.205 -48.05 9.295 -47.042 ;
      RECT 9.155 -47.815 9.295 -47.645 ;
      RECT 9.205 -46.628 9.295 -45.62 ;
      RECT 9.155 -46.025 9.295 -45.855 ;
      RECT 9.205 -44.82 9.295 -43.812 ;
      RECT 9.155 -44.585 9.295 -44.415 ;
      RECT 9.205 -43.398 9.295 -42.39 ;
      RECT 9.155 -42.795 9.295 -42.625 ;
      RECT 9.205 -41.59 9.295 -40.582 ;
      RECT 9.155 -41.355 9.295 -41.185 ;
      RECT 9.205 -40.168 9.295 -39.16 ;
      RECT 9.155 -39.565 9.295 -39.395 ;
      RECT 9.205 -38.36 9.295 -37.352 ;
      RECT 9.155 -38.125 9.295 -37.955 ;
      RECT 9.205 -36.938 9.295 -35.93 ;
      RECT 9.155 -36.335 9.295 -36.165 ;
      RECT 9.205 -35.13 9.295 -34.122 ;
      RECT 9.155 -34.895 9.295 -34.725 ;
      RECT 9.205 -33.708 9.295 -32.7 ;
      RECT 9.155 -33.105 9.295 -32.935 ;
      RECT 9.205 -31.9 9.295 -30.892 ;
      RECT 9.155 -31.665 9.295 -31.495 ;
      RECT 9.205 -30.478 9.295 -29.47 ;
      RECT 9.155 -29.875 9.295 -29.705 ;
      RECT 9.205 -28.67 9.295 -27.662 ;
      RECT 9.155 -28.435 9.295 -28.265 ;
      RECT 9.205 -27.248 9.295 -26.24 ;
      RECT 9.155 -26.645 9.295 -26.475 ;
      RECT 9.205 -25.44 9.295 -24.432 ;
      RECT 9.155 -25.205 9.295 -25.035 ;
      RECT 9.205 -24.018 9.295 -23.01 ;
      RECT 9.155 -23.415 9.295 -23.245 ;
      RECT 9.205 -22.21 9.295 -21.202 ;
      RECT 9.155 -21.975 9.295 -21.805 ;
      RECT 9.205 -20.788 9.295 -19.78 ;
      RECT 9.155 -20.185 9.295 -20.015 ;
      RECT 9.205 -18.98 9.295 -17.972 ;
      RECT 9.155 -18.745 9.295 -18.575 ;
      RECT 9.205 -17.558 9.295 -16.55 ;
      RECT 9.155 -16.955 9.295 -16.785 ;
      RECT 9.205 -15.75 9.295 -14.742 ;
      RECT 9.155 -15.515 9.295 -15.345 ;
      RECT 9.205 -14.328 9.295 -13.32 ;
      RECT 9.155 -13.725 9.295 -13.555 ;
      RECT 9.205 -12.52 9.295 -11.512 ;
      RECT 9.155 -12.285 9.295 -12.115 ;
      RECT 9.205 -11.098 9.295 -10.09 ;
      RECT 9.155 -10.495 9.295 -10.325 ;
      RECT 9.205 -9.29 9.295 -8.282 ;
      RECT 9.155 -9.055 9.295 -8.885 ;
      RECT 9.205 -7.868 9.295 -6.86 ;
      RECT 9.155 -7.265 9.295 -7.095 ;
      RECT 9.205 -6.06 9.295 -5.052 ;
      RECT 9.155 -5.825 9.295 -5.655 ;
      RECT 9.205 -4.638 9.295 -3.63 ;
      RECT 9.155 -4.035 9.295 -3.865 ;
      RECT 9.205 -2.83 9.295 -1.822 ;
      RECT 9.155 -2.595 9.295 -2.425 ;
      RECT 9.205 -1.408 9.295 -0.4 ;
      RECT 9.155 -0.805 9.295 -0.635 ;
      RECT 9.205 0.4 9.295 1.408 ;
      RECT 9.155 0.635 9.295 0.805 ;
      RECT 7.775 -60.005 9.255 -59.905 ;
      RECT 7.775 -60.515 7.875 -59.905 ;
      RECT 7.995 -57.47 9.255 -57.37 ;
      RECT 9.155 -57.795 9.255 -57.37 ;
      RECT 8.595 -57.795 8.695 -57.37 ;
      RECT 8.035 -57.795 8.135 -57.37 ;
      RECT 8.805 -49.858 8.895 -48.851 ;
      RECT 8.805 -49.545 8.945 -49.375 ;
      RECT 8.805 -48.049 8.895 -47.042 ;
      RECT 8.805 -47.525 8.945 -47.355 ;
      RECT 8.805 -46.628 8.895 -45.621 ;
      RECT 8.805 -46.315 8.945 -46.145 ;
      RECT 8.805 -44.819 8.895 -43.812 ;
      RECT 8.805 -44.295 8.945 -44.125 ;
      RECT 8.805 -43.398 8.895 -42.391 ;
      RECT 8.805 -43.085 8.945 -42.915 ;
      RECT 8.805 -41.589 8.895 -40.582 ;
      RECT 8.805 -41.065 8.945 -40.895 ;
      RECT 8.805 -40.168 8.895 -39.161 ;
      RECT 8.805 -39.855 8.945 -39.685 ;
      RECT 8.805 -38.359 8.895 -37.352 ;
      RECT 8.805 -37.835 8.945 -37.665 ;
      RECT 8.805 -36.938 8.895 -35.931 ;
      RECT 8.805 -36.625 8.945 -36.455 ;
      RECT 8.805 -35.129 8.895 -34.122 ;
      RECT 8.805 -34.605 8.945 -34.435 ;
      RECT 8.805 -33.708 8.895 -32.701 ;
      RECT 8.805 -33.395 8.945 -33.225 ;
      RECT 8.805 -31.899 8.895 -30.892 ;
      RECT 8.805 -31.375 8.945 -31.205 ;
      RECT 8.805 -30.478 8.895 -29.471 ;
      RECT 8.805 -30.165 8.945 -29.995 ;
      RECT 8.805 -28.669 8.895 -27.662 ;
      RECT 8.805 -28.145 8.945 -27.975 ;
      RECT 8.805 -27.248 8.895 -26.241 ;
      RECT 8.805 -26.935 8.945 -26.765 ;
      RECT 8.805 -25.439 8.895 -24.432 ;
      RECT 8.805 -24.915 8.945 -24.745 ;
      RECT 8.805 -24.018 8.895 -23.011 ;
      RECT 8.805 -23.705 8.945 -23.535 ;
      RECT 8.805 -22.209 8.895 -21.202 ;
      RECT 8.805 -21.685 8.945 -21.515 ;
      RECT 8.805 -20.788 8.895 -19.781 ;
      RECT 8.805 -20.475 8.945 -20.305 ;
      RECT 8.805 -18.979 8.895 -17.972 ;
      RECT 8.805 -18.455 8.945 -18.285 ;
      RECT 8.805 -17.558 8.895 -16.551 ;
      RECT 8.805 -17.245 8.945 -17.075 ;
      RECT 8.805 -15.749 8.895 -14.742 ;
      RECT 8.805 -15.225 8.945 -15.055 ;
      RECT 8.805 -14.328 8.895 -13.321 ;
      RECT 8.805 -14.015 8.945 -13.845 ;
      RECT 8.805 -12.519 8.895 -11.512 ;
      RECT 8.805 -11.995 8.945 -11.825 ;
      RECT 8.805 -11.098 8.895 -10.091 ;
      RECT 8.805 -10.785 8.945 -10.615 ;
      RECT 8.805 -9.289 8.895 -8.282 ;
      RECT 8.805 -8.765 8.945 -8.595 ;
      RECT 8.805 -7.868 8.895 -6.861 ;
      RECT 8.805 -7.555 8.945 -7.385 ;
      RECT 8.805 -6.059 8.895 -5.052 ;
      RECT 8.805 -5.535 8.945 -5.365 ;
      RECT 8.805 -4.638 8.895 -3.631 ;
      RECT 8.805 -4.325 8.945 -4.155 ;
      RECT 8.805 -2.829 8.895 -1.822 ;
      RECT 8.805 -2.305 8.945 -2.135 ;
      RECT 8.805 -1.408 8.895 -0.401 ;
      RECT 8.805 -1.095 8.945 -0.925 ;
      RECT 8.805 0.401 8.895 1.408 ;
      RECT 8.805 0.925 8.945 1.095 ;
      RECT 8.135 -59.815 8.305 -59.705 ;
      RECT 4.985 -59.815 8.305 -59.715 ;
      RECT 8.005 -49.858 8.095 -48.85 ;
      RECT 7.955 -49.255 8.095 -49.085 ;
      RECT 8.005 -48.05 8.095 -47.042 ;
      RECT 7.955 -47.815 8.095 -47.645 ;
      RECT 8.005 -46.628 8.095 -45.62 ;
      RECT 7.955 -46.025 8.095 -45.855 ;
      RECT 8.005 -44.82 8.095 -43.812 ;
      RECT 7.955 -44.585 8.095 -44.415 ;
      RECT 8.005 -43.398 8.095 -42.39 ;
      RECT 7.955 -42.795 8.095 -42.625 ;
      RECT 8.005 -41.59 8.095 -40.582 ;
      RECT 7.955 -41.355 8.095 -41.185 ;
      RECT 8.005 -40.168 8.095 -39.16 ;
      RECT 7.955 -39.565 8.095 -39.395 ;
      RECT 8.005 -38.36 8.095 -37.352 ;
      RECT 7.955 -38.125 8.095 -37.955 ;
      RECT 8.005 -36.938 8.095 -35.93 ;
      RECT 7.955 -36.335 8.095 -36.165 ;
      RECT 8.005 -35.13 8.095 -34.122 ;
      RECT 7.955 -34.895 8.095 -34.725 ;
      RECT 8.005 -33.708 8.095 -32.7 ;
      RECT 7.955 -33.105 8.095 -32.935 ;
      RECT 8.005 -31.9 8.095 -30.892 ;
      RECT 7.955 -31.665 8.095 -31.495 ;
      RECT 8.005 -30.478 8.095 -29.47 ;
      RECT 7.955 -29.875 8.095 -29.705 ;
      RECT 8.005 -28.67 8.095 -27.662 ;
      RECT 7.955 -28.435 8.095 -28.265 ;
      RECT 8.005 -27.248 8.095 -26.24 ;
      RECT 7.955 -26.645 8.095 -26.475 ;
      RECT 8.005 -25.44 8.095 -24.432 ;
      RECT 7.955 -25.205 8.095 -25.035 ;
      RECT 8.005 -24.018 8.095 -23.01 ;
      RECT 7.955 -23.415 8.095 -23.245 ;
      RECT 8.005 -22.21 8.095 -21.202 ;
      RECT 7.955 -21.975 8.095 -21.805 ;
      RECT 8.005 -20.788 8.095 -19.78 ;
      RECT 7.955 -20.185 8.095 -20.015 ;
      RECT 8.005 -18.98 8.095 -17.972 ;
      RECT 7.955 -18.745 8.095 -18.575 ;
      RECT 8.005 -17.558 8.095 -16.55 ;
      RECT 7.955 -16.955 8.095 -16.785 ;
      RECT 8.005 -15.75 8.095 -14.742 ;
      RECT 7.955 -15.515 8.095 -15.345 ;
      RECT 8.005 -14.328 8.095 -13.32 ;
      RECT 7.955 -13.725 8.095 -13.555 ;
      RECT 8.005 -12.52 8.095 -11.512 ;
      RECT 7.955 -12.285 8.095 -12.115 ;
      RECT 8.005 -11.098 8.095 -10.09 ;
      RECT 7.955 -10.495 8.095 -10.325 ;
      RECT 8.005 -9.29 8.095 -8.282 ;
      RECT 7.955 -9.055 8.095 -8.885 ;
      RECT 8.005 -7.868 8.095 -6.86 ;
      RECT 7.955 -7.265 8.095 -7.095 ;
      RECT 8.005 -6.06 8.095 -5.052 ;
      RECT 7.955 -5.825 8.095 -5.655 ;
      RECT 8.005 -4.638 8.095 -3.63 ;
      RECT 7.955 -4.035 8.095 -3.865 ;
      RECT 8.005 -2.83 8.095 -1.822 ;
      RECT 7.955 -2.595 8.095 -2.425 ;
      RECT 8.005 -1.408 8.095 -0.4 ;
      RECT 7.955 -0.805 8.095 -0.635 ;
      RECT 8.005 0.4 8.095 1.408 ;
      RECT 7.955 0.635 8.095 0.805 ;
      RECT 7.605 -49.858 7.695 -48.851 ;
      RECT 7.605 -49.545 7.745 -49.375 ;
      RECT 7.605 -48.049 7.695 -47.042 ;
      RECT 7.605 -47.525 7.745 -47.355 ;
      RECT 7.605 -46.628 7.695 -45.621 ;
      RECT 7.605 -46.315 7.745 -46.145 ;
      RECT 7.605 -44.819 7.695 -43.812 ;
      RECT 7.605 -44.295 7.745 -44.125 ;
      RECT 7.605 -43.398 7.695 -42.391 ;
      RECT 7.605 -43.085 7.745 -42.915 ;
      RECT 7.605 -41.589 7.695 -40.582 ;
      RECT 7.605 -41.065 7.745 -40.895 ;
      RECT 7.605 -40.168 7.695 -39.161 ;
      RECT 7.605 -39.855 7.745 -39.685 ;
      RECT 7.605 -38.359 7.695 -37.352 ;
      RECT 7.605 -37.835 7.745 -37.665 ;
      RECT 7.605 -36.938 7.695 -35.931 ;
      RECT 7.605 -36.625 7.745 -36.455 ;
      RECT 7.605 -35.129 7.695 -34.122 ;
      RECT 7.605 -34.605 7.745 -34.435 ;
      RECT 7.605 -33.708 7.695 -32.701 ;
      RECT 7.605 -33.395 7.745 -33.225 ;
      RECT 7.605 -31.899 7.695 -30.892 ;
      RECT 7.605 -31.375 7.745 -31.205 ;
      RECT 7.605 -30.478 7.695 -29.471 ;
      RECT 7.605 -30.165 7.745 -29.995 ;
      RECT 7.605 -28.669 7.695 -27.662 ;
      RECT 7.605 -28.145 7.745 -27.975 ;
      RECT 7.605 -27.248 7.695 -26.241 ;
      RECT 7.605 -26.935 7.745 -26.765 ;
      RECT 7.605 -25.439 7.695 -24.432 ;
      RECT 7.605 -24.915 7.745 -24.745 ;
      RECT 7.605 -24.018 7.695 -23.011 ;
      RECT 7.605 -23.705 7.745 -23.535 ;
      RECT 7.605 -22.209 7.695 -21.202 ;
      RECT 7.605 -21.685 7.745 -21.515 ;
      RECT 7.605 -20.788 7.695 -19.781 ;
      RECT 7.605 -20.475 7.745 -20.305 ;
      RECT 7.605 -18.979 7.695 -17.972 ;
      RECT 7.605 -18.455 7.745 -18.285 ;
      RECT 7.605 -17.558 7.695 -16.551 ;
      RECT 7.605 -17.245 7.745 -17.075 ;
      RECT 7.605 -15.749 7.695 -14.742 ;
      RECT 7.605 -15.225 7.745 -15.055 ;
      RECT 7.605 -14.328 7.695 -13.321 ;
      RECT 7.605 -14.015 7.745 -13.845 ;
      RECT 7.605 -12.519 7.695 -11.512 ;
      RECT 7.605 -11.995 7.745 -11.825 ;
      RECT 7.605 -11.098 7.695 -10.091 ;
      RECT 7.605 -10.785 7.745 -10.615 ;
      RECT 7.605 -9.289 7.695 -8.282 ;
      RECT 7.605 -8.765 7.745 -8.595 ;
      RECT 7.605 -7.868 7.695 -6.861 ;
      RECT 7.605 -7.555 7.745 -7.385 ;
      RECT 7.605 -6.059 7.695 -5.052 ;
      RECT 7.605 -5.535 7.745 -5.365 ;
      RECT 7.605 -4.638 7.695 -3.631 ;
      RECT 7.605 -4.325 7.745 -4.155 ;
      RECT 7.605 -2.829 7.695 -1.822 ;
      RECT 7.605 -2.305 7.745 -2.135 ;
      RECT 7.605 -1.408 7.695 -0.401 ;
      RECT 7.605 -1.095 7.745 -0.925 ;
      RECT 7.605 0.401 7.695 1.408 ;
      RECT 7.605 0.925 7.745 1.095 ;
      RECT 5.755 -60.005 7.235 -59.905 ;
      RECT 5.755 -60.375 5.855 -59.905 ;
      RECT 5.56 -62.715 7.135 -62.595 ;
      RECT 7.035 -63.215 7.135 -62.595 ;
      RECT 6.44 -63.215 6.54 -62.595 ;
      RECT 5.56 -63.17 5.66 -62.595 ;
      RECT 6.805 -49.858 6.895 -48.85 ;
      RECT 6.755 -49.255 6.895 -49.085 ;
      RECT 6.805 -48.05 6.895 -47.042 ;
      RECT 6.755 -47.815 6.895 -47.645 ;
      RECT 6.805 -46.628 6.895 -45.62 ;
      RECT 6.755 -46.025 6.895 -45.855 ;
      RECT 6.805 -44.82 6.895 -43.812 ;
      RECT 6.755 -44.585 6.895 -44.415 ;
      RECT 6.805 -43.398 6.895 -42.39 ;
      RECT 6.755 -42.795 6.895 -42.625 ;
      RECT 6.805 -41.59 6.895 -40.582 ;
      RECT 6.755 -41.355 6.895 -41.185 ;
      RECT 6.805 -40.168 6.895 -39.16 ;
      RECT 6.755 -39.565 6.895 -39.395 ;
      RECT 6.805 -38.36 6.895 -37.352 ;
      RECT 6.755 -38.125 6.895 -37.955 ;
      RECT 6.805 -36.938 6.895 -35.93 ;
      RECT 6.755 -36.335 6.895 -36.165 ;
      RECT 6.805 -35.13 6.895 -34.122 ;
      RECT 6.755 -34.895 6.895 -34.725 ;
      RECT 6.805 -33.708 6.895 -32.7 ;
      RECT 6.755 -33.105 6.895 -32.935 ;
      RECT 6.805 -31.9 6.895 -30.892 ;
      RECT 6.755 -31.665 6.895 -31.495 ;
      RECT 6.805 -30.478 6.895 -29.47 ;
      RECT 6.755 -29.875 6.895 -29.705 ;
      RECT 6.805 -28.67 6.895 -27.662 ;
      RECT 6.755 -28.435 6.895 -28.265 ;
      RECT 6.805 -27.248 6.895 -26.24 ;
      RECT 6.755 -26.645 6.895 -26.475 ;
      RECT 6.805 -25.44 6.895 -24.432 ;
      RECT 6.755 -25.205 6.895 -25.035 ;
      RECT 6.805 -24.018 6.895 -23.01 ;
      RECT 6.755 -23.415 6.895 -23.245 ;
      RECT 6.805 -22.21 6.895 -21.202 ;
      RECT 6.755 -21.975 6.895 -21.805 ;
      RECT 6.805 -20.788 6.895 -19.78 ;
      RECT 6.755 -20.185 6.895 -20.015 ;
      RECT 6.805 -18.98 6.895 -17.972 ;
      RECT 6.755 -18.745 6.895 -18.575 ;
      RECT 6.805 -17.558 6.895 -16.55 ;
      RECT 6.755 -16.955 6.895 -16.785 ;
      RECT 6.805 -15.75 6.895 -14.742 ;
      RECT 6.755 -15.515 6.895 -15.345 ;
      RECT 6.805 -14.328 6.895 -13.32 ;
      RECT 6.755 -13.725 6.895 -13.555 ;
      RECT 6.805 -12.52 6.895 -11.512 ;
      RECT 6.755 -12.285 6.895 -12.115 ;
      RECT 6.805 -11.098 6.895 -10.09 ;
      RECT 6.755 -10.495 6.895 -10.325 ;
      RECT 6.805 -9.29 6.895 -8.282 ;
      RECT 6.755 -9.055 6.895 -8.885 ;
      RECT 6.805 -7.868 6.895 -6.86 ;
      RECT 6.755 -7.265 6.895 -7.095 ;
      RECT 6.805 -6.06 6.895 -5.052 ;
      RECT 6.755 -5.825 6.895 -5.655 ;
      RECT 6.805 -4.638 6.895 -3.63 ;
      RECT 6.755 -4.035 6.895 -3.865 ;
      RECT 6.805 -2.83 6.895 -1.822 ;
      RECT 6.755 -2.595 6.895 -2.425 ;
      RECT 6.805 -1.408 6.895 -0.4 ;
      RECT 6.755 -0.805 6.895 -0.635 ;
      RECT 6.805 0.4 6.895 1.408 ;
      RECT 6.755 0.635 6.895 0.805 ;
      RECT 6.68 -63.005 6.855 -62.835 ;
      RECT 6.755 -63.215 6.855 -62.835 ;
      RECT 5.795 -61.875 5.895 -61.41 ;
      RECT 6.16 -61.875 6.26 -61.42 ;
      RECT 5.795 -61.875 6.64 -61.705 ;
      RECT 6.405 -49.858 6.495 -48.851 ;
      RECT 6.405 -49.545 6.545 -49.375 ;
      RECT 6.405 -48.049 6.495 -47.042 ;
      RECT 6.405 -47.525 6.545 -47.355 ;
      RECT 6.405 -46.628 6.495 -45.621 ;
      RECT 6.405 -46.315 6.545 -46.145 ;
      RECT 6.405 -44.819 6.495 -43.812 ;
      RECT 6.405 -44.295 6.545 -44.125 ;
      RECT 6.405 -43.398 6.495 -42.391 ;
      RECT 6.405 -43.085 6.545 -42.915 ;
      RECT 6.405 -41.589 6.495 -40.582 ;
      RECT 6.405 -41.065 6.545 -40.895 ;
      RECT 6.405 -40.168 6.495 -39.161 ;
      RECT 6.405 -39.855 6.545 -39.685 ;
      RECT 6.405 -38.359 6.495 -37.352 ;
      RECT 6.405 -37.835 6.545 -37.665 ;
      RECT 6.405 -36.938 6.495 -35.931 ;
      RECT 6.405 -36.625 6.545 -36.455 ;
      RECT 6.405 -35.129 6.495 -34.122 ;
      RECT 6.405 -34.605 6.545 -34.435 ;
      RECT 6.405 -33.708 6.495 -32.701 ;
      RECT 6.405 -33.395 6.545 -33.225 ;
      RECT 6.405 -31.899 6.495 -30.892 ;
      RECT 6.405 -31.375 6.545 -31.205 ;
      RECT 6.405 -30.478 6.495 -29.471 ;
      RECT 6.405 -30.165 6.545 -29.995 ;
      RECT 6.405 -28.669 6.495 -27.662 ;
      RECT 6.405 -28.145 6.545 -27.975 ;
      RECT 6.405 -27.248 6.495 -26.241 ;
      RECT 6.405 -26.935 6.545 -26.765 ;
      RECT 6.405 -25.439 6.495 -24.432 ;
      RECT 6.405 -24.915 6.545 -24.745 ;
      RECT 6.405 -24.018 6.495 -23.011 ;
      RECT 6.405 -23.705 6.545 -23.535 ;
      RECT 6.405 -22.209 6.495 -21.202 ;
      RECT 6.405 -21.685 6.545 -21.515 ;
      RECT 6.405 -20.788 6.495 -19.781 ;
      RECT 6.405 -20.475 6.545 -20.305 ;
      RECT 6.405 -18.979 6.495 -17.972 ;
      RECT 6.405 -18.455 6.545 -18.285 ;
      RECT 6.405 -17.558 6.495 -16.551 ;
      RECT 6.405 -17.245 6.545 -17.075 ;
      RECT 6.405 -15.749 6.495 -14.742 ;
      RECT 6.405 -15.225 6.545 -15.055 ;
      RECT 6.405 -14.328 6.495 -13.321 ;
      RECT 6.405 -14.015 6.545 -13.845 ;
      RECT 6.405 -12.519 6.495 -11.512 ;
      RECT 6.405 -11.995 6.545 -11.825 ;
      RECT 6.405 -11.098 6.495 -10.091 ;
      RECT 6.405 -10.785 6.545 -10.615 ;
      RECT 6.405 -9.289 6.495 -8.282 ;
      RECT 6.405 -8.765 6.545 -8.595 ;
      RECT 6.405 -7.868 6.495 -6.861 ;
      RECT 6.405 -7.555 6.545 -7.385 ;
      RECT 6.405 -6.059 6.495 -5.052 ;
      RECT 6.405 -5.535 6.545 -5.365 ;
      RECT 6.405 -4.638 6.495 -3.631 ;
      RECT 6.405 -4.325 6.545 -4.155 ;
      RECT 6.405 -2.829 6.495 -1.822 ;
      RECT 6.405 -2.305 6.545 -2.135 ;
      RECT 6.405 -1.408 6.495 -0.401 ;
      RECT 6.405 -1.095 6.545 -0.925 ;
      RECT 6.405 0.401 6.495 1.408 ;
      RECT 6.405 0.925 6.545 1.095 ;
      RECT 6.09 -63.005 6.26 -62.835 ;
      RECT 6.16 -63.215 6.26 -62.835 ;
      RECT 5.605 -49.858 5.695 -48.85 ;
      RECT 5.555 -49.255 5.695 -49.085 ;
      RECT 5.605 -48.05 5.695 -47.042 ;
      RECT 5.555 -47.815 5.695 -47.645 ;
      RECT 5.605 -46.628 5.695 -45.62 ;
      RECT 5.555 -46.025 5.695 -45.855 ;
      RECT 5.605 -44.82 5.695 -43.812 ;
      RECT 5.555 -44.585 5.695 -44.415 ;
      RECT 5.605 -43.398 5.695 -42.39 ;
      RECT 5.555 -42.795 5.695 -42.625 ;
      RECT 5.605 -41.59 5.695 -40.582 ;
      RECT 5.555 -41.355 5.695 -41.185 ;
      RECT 5.605 -40.168 5.695 -39.16 ;
      RECT 5.555 -39.565 5.695 -39.395 ;
      RECT 5.605 -38.36 5.695 -37.352 ;
      RECT 5.555 -38.125 5.695 -37.955 ;
      RECT 5.605 -36.938 5.695 -35.93 ;
      RECT 5.555 -36.335 5.695 -36.165 ;
      RECT 5.605 -35.13 5.695 -34.122 ;
      RECT 5.555 -34.895 5.695 -34.725 ;
      RECT 5.605 -33.708 5.695 -32.7 ;
      RECT 5.555 -33.105 5.695 -32.935 ;
      RECT 5.605 -31.9 5.695 -30.892 ;
      RECT 5.555 -31.665 5.695 -31.495 ;
      RECT 5.605 -30.478 5.695 -29.47 ;
      RECT 5.555 -29.875 5.695 -29.705 ;
      RECT 5.605 -28.67 5.695 -27.662 ;
      RECT 5.555 -28.435 5.695 -28.265 ;
      RECT 5.605 -27.248 5.695 -26.24 ;
      RECT 5.555 -26.645 5.695 -26.475 ;
      RECT 5.605 -25.44 5.695 -24.432 ;
      RECT 5.555 -25.205 5.695 -25.035 ;
      RECT 5.605 -24.018 5.695 -23.01 ;
      RECT 5.555 -23.415 5.695 -23.245 ;
      RECT 5.605 -22.21 5.695 -21.202 ;
      RECT 5.555 -21.975 5.695 -21.805 ;
      RECT 5.605 -20.788 5.695 -19.78 ;
      RECT 5.555 -20.185 5.695 -20.015 ;
      RECT 5.605 -18.98 5.695 -17.972 ;
      RECT 5.555 -18.745 5.695 -18.575 ;
      RECT 5.605 -17.558 5.695 -16.55 ;
      RECT 5.555 -16.955 5.695 -16.785 ;
      RECT 5.605 -15.75 5.695 -14.742 ;
      RECT 5.555 -15.515 5.695 -15.345 ;
      RECT 5.605 -14.328 5.695 -13.32 ;
      RECT 5.555 -13.725 5.695 -13.555 ;
      RECT 5.605 -12.52 5.695 -11.512 ;
      RECT 5.555 -12.285 5.695 -12.115 ;
      RECT 5.605 -11.098 5.695 -10.09 ;
      RECT 5.555 -10.495 5.695 -10.325 ;
      RECT 5.605 -9.29 5.695 -8.282 ;
      RECT 5.555 -9.055 5.695 -8.885 ;
      RECT 5.605 -7.868 5.695 -6.86 ;
      RECT 5.555 -7.265 5.695 -7.095 ;
      RECT 5.605 -6.06 5.695 -5.052 ;
      RECT 5.555 -5.825 5.695 -5.655 ;
      RECT 5.605 -4.638 5.695 -3.63 ;
      RECT 5.555 -4.035 5.695 -3.865 ;
      RECT 5.605 -2.83 5.695 -1.822 ;
      RECT 5.555 -2.595 5.695 -2.425 ;
      RECT 5.605 -1.408 5.695 -0.4 ;
      RECT 5.555 -0.805 5.695 -0.635 ;
      RECT 5.605 0.4 5.695 1.408 ;
      RECT 5.555 0.635 5.695 0.805 ;
      RECT 5.205 -49.858 5.295 -48.851 ;
      RECT 5.205 -49.545 5.345 -49.375 ;
      RECT 5.205 -48.049 5.295 -47.042 ;
      RECT 5.205 -47.525 5.345 -47.355 ;
      RECT 5.205 -46.628 5.295 -45.621 ;
      RECT 5.205 -46.315 5.345 -46.145 ;
      RECT 5.205 -44.819 5.295 -43.812 ;
      RECT 5.205 -44.295 5.345 -44.125 ;
      RECT 5.205 -43.398 5.295 -42.391 ;
      RECT 5.205 -43.085 5.345 -42.915 ;
      RECT 5.205 -41.589 5.295 -40.582 ;
      RECT 5.205 -41.065 5.345 -40.895 ;
      RECT 5.205 -40.168 5.295 -39.161 ;
      RECT 5.205 -39.855 5.345 -39.685 ;
      RECT 5.205 -38.359 5.295 -37.352 ;
      RECT 5.205 -37.835 5.345 -37.665 ;
      RECT 5.205 -36.938 5.295 -35.931 ;
      RECT 5.205 -36.625 5.345 -36.455 ;
      RECT 5.205 -35.129 5.295 -34.122 ;
      RECT 5.205 -34.605 5.345 -34.435 ;
      RECT 5.205 -33.708 5.295 -32.701 ;
      RECT 5.205 -33.395 5.345 -33.225 ;
      RECT 5.205 -31.899 5.295 -30.892 ;
      RECT 5.205 -31.375 5.345 -31.205 ;
      RECT 5.205 -30.478 5.295 -29.471 ;
      RECT 5.205 -30.165 5.345 -29.995 ;
      RECT 5.205 -28.669 5.295 -27.662 ;
      RECT 5.205 -28.145 5.345 -27.975 ;
      RECT 5.205 -27.248 5.295 -26.241 ;
      RECT 5.205 -26.935 5.345 -26.765 ;
      RECT 5.205 -25.439 5.295 -24.432 ;
      RECT 5.205 -24.915 5.345 -24.745 ;
      RECT 5.205 -24.018 5.295 -23.011 ;
      RECT 5.205 -23.705 5.345 -23.535 ;
      RECT 5.205 -22.209 5.295 -21.202 ;
      RECT 5.205 -21.685 5.345 -21.515 ;
      RECT 5.205 -20.788 5.295 -19.781 ;
      RECT 5.205 -20.475 5.345 -20.305 ;
      RECT 5.205 -18.979 5.295 -17.972 ;
      RECT 5.205 -18.455 5.345 -18.285 ;
      RECT 5.205 -17.558 5.295 -16.551 ;
      RECT 5.205 -17.245 5.345 -17.075 ;
      RECT 5.205 -15.749 5.295 -14.742 ;
      RECT 5.205 -15.225 5.345 -15.055 ;
      RECT 5.205 -14.328 5.295 -13.321 ;
      RECT 5.205 -14.015 5.345 -13.845 ;
      RECT 5.205 -12.519 5.295 -11.512 ;
      RECT 5.205 -11.995 5.345 -11.825 ;
      RECT 5.205 -11.098 5.295 -10.091 ;
      RECT 5.205 -10.785 5.345 -10.615 ;
      RECT 5.205 -9.289 5.295 -8.282 ;
      RECT 5.205 -8.765 5.345 -8.595 ;
      RECT 5.205 -7.868 5.295 -6.861 ;
      RECT 5.205 -7.555 5.345 -7.385 ;
      RECT 5.205 -6.059 5.295 -5.052 ;
      RECT 5.205 -5.535 5.345 -5.365 ;
      RECT 5.205 -4.638 5.295 -3.631 ;
      RECT 5.205 -4.325 5.345 -4.155 ;
      RECT 5.205 -2.829 5.295 -1.822 ;
      RECT 5.205 -2.305 5.345 -2.135 ;
      RECT 5.205 -1.408 5.295 -0.401 ;
      RECT 5.205 -1.095 5.345 -0.925 ;
      RECT 5.205 0.401 5.295 1.408 ;
      RECT 5.205 0.925 5.345 1.095 ;
      RECT 1.035 -57.255 4.815 -57.135 ;
      RECT 2.355 -57.795 2.455 -57.135 ;
      RECT 1.795 -57.795 1.895 -57.135 ;
      RECT 1.235 -57.795 1.335 -57.135 ;
      RECT 4.405 -49.858 4.495 -48.85 ;
      RECT 4.355 -49.255 4.495 -49.085 ;
      RECT 4.405 -48.05 4.495 -47.042 ;
      RECT 4.355 -47.815 4.495 -47.645 ;
      RECT 4.405 -46.628 4.495 -45.62 ;
      RECT 4.355 -46.025 4.495 -45.855 ;
      RECT 4.405 -44.82 4.495 -43.812 ;
      RECT 4.355 -44.585 4.495 -44.415 ;
      RECT 4.405 -43.398 4.495 -42.39 ;
      RECT 4.355 -42.795 4.495 -42.625 ;
      RECT 4.405 -41.59 4.495 -40.582 ;
      RECT 4.355 -41.355 4.495 -41.185 ;
      RECT 4.405 -40.168 4.495 -39.16 ;
      RECT 4.355 -39.565 4.495 -39.395 ;
      RECT 4.405 -38.36 4.495 -37.352 ;
      RECT 4.355 -38.125 4.495 -37.955 ;
      RECT 4.405 -36.938 4.495 -35.93 ;
      RECT 4.355 -36.335 4.495 -36.165 ;
      RECT 4.405 -35.13 4.495 -34.122 ;
      RECT 4.355 -34.895 4.495 -34.725 ;
      RECT 4.405 -33.708 4.495 -32.7 ;
      RECT 4.355 -33.105 4.495 -32.935 ;
      RECT 4.405 -31.9 4.495 -30.892 ;
      RECT 4.355 -31.665 4.495 -31.495 ;
      RECT 4.405 -30.478 4.495 -29.47 ;
      RECT 4.355 -29.875 4.495 -29.705 ;
      RECT 4.405 -28.67 4.495 -27.662 ;
      RECT 4.355 -28.435 4.495 -28.265 ;
      RECT 4.405 -27.248 4.495 -26.24 ;
      RECT 4.355 -26.645 4.495 -26.475 ;
      RECT 4.405 -25.44 4.495 -24.432 ;
      RECT 4.355 -25.205 4.495 -25.035 ;
      RECT 4.405 -24.018 4.495 -23.01 ;
      RECT 4.355 -23.415 4.495 -23.245 ;
      RECT 4.405 -22.21 4.495 -21.202 ;
      RECT 4.355 -21.975 4.495 -21.805 ;
      RECT 4.405 -20.788 4.495 -19.78 ;
      RECT 4.355 -20.185 4.495 -20.015 ;
      RECT 4.405 -18.98 4.495 -17.972 ;
      RECT 4.355 -18.745 4.495 -18.575 ;
      RECT 4.405 -17.558 4.495 -16.55 ;
      RECT 4.355 -16.955 4.495 -16.785 ;
      RECT 4.405 -15.75 4.495 -14.742 ;
      RECT 4.355 -15.515 4.495 -15.345 ;
      RECT 4.405 -14.328 4.495 -13.32 ;
      RECT 4.355 -13.725 4.495 -13.555 ;
      RECT 4.405 -12.52 4.495 -11.512 ;
      RECT 4.355 -12.285 4.495 -12.115 ;
      RECT 4.405 -11.098 4.495 -10.09 ;
      RECT 4.355 -10.495 4.495 -10.325 ;
      RECT 4.405 -9.29 4.495 -8.282 ;
      RECT 4.355 -9.055 4.495 -8.885 ;
      RECT 4.405 -7.868 4.495 -6.86 ;
      RECT 4.355 -7.265 4.495 -7.095 ;
      RECT 4.405 -6.06 4.495 -5.052 ;
      RECT 4.355 -5.825 4.495 -5.655 ;
      RECT 4.405 -4.638 4.495 -3.63 ;
      RECT 4.355 -4.035 4.495 -3.865 ;
      RECT 4.405 -2.83 4.495 -1.822 ;
      RECT 4.355 -2.595 4.495 -2.425 ;
      RECT 4.405 -1.408 4.495 -0.4 ;
      RECT 4.355 -0.805 4.495 -0.635 ;
      RECT 4.405 0.4 4.495 1.408 ;
      RECT 4.355 0.635 4.495 0.805 ;
      RECT 2.975 -60.005 4.455 -59.905 ;
      RECT 2.975 -60.515 3.075 -59.905 ;
      RECT 3.195 -57.47 4.455 -57.37 ;
      RECT 4.355 -57.795 4.455 -57.37 ;
      RECT 3.795 -57.795 3.895 -57.37 ;
      RECT 3.235 -57.795 3.335 -57.37 ;
      RECT 4.005 -49.858 4.095 -48.851 ;
      RECT 4.005 -49.545 4.145 -49.375 ;
      RECT 4.005 -48.049 4.095 -47.042 ;
      RECT 4.005 -47.525 4.145 -47.355 ;
      RECT 4.005 -46.628 4.095 -45.621 ;
      RECT 4.005 -46.315 4.145 -46.145 ;
      RECT 4.005 -44.819 4.095 -43.812 ;
      RECT 4.005 -44.295 4.145 -44.125 ;
      RECT 4.005 -43.398 4.095 -42.391 ;
      RECT 4.005 -43.085 4.145 -42.915 ;
      RECT 4.005 -41.589 4.095 -40.582 ;
      RECT 4.005 -41.065 4.145 -40.895 ;
      RECT 4.005 -40.168 4.095 -39.161 ;
      RECT 4.005 -39.855 4.145 -39.685 ;
      RECT 4.005 -38.359 4.095 -37.352 ;
      RECT 4.005 -37.835 4.145 -37.665 ;
      RECT 4.005 -36.938 4.095 -35.931 ;
      RECT 4.005 -36.625 4.145 -36.455 ;
      RECT 4.005 -35.129 4.095 -34.122 ;
      RECT 4.005 -34.605 4.145 -34.435 ;
      RECT 4.005 -33.708 4.095 -32.701 ;
      RECT 4.005 -33.395 4.145 -33.225 ;
      RECT 4.005 -31.899 4.095 -30.892 ;
      RECT 4.005 -31.375 4.145 -31.205 ;
      RECT 4.005 -30.478 4.095 -29.471 ;
      RECT 4.005 -30.165 4.145 -29.995 ;
      RECT 4.005 -28.669 4.095 -27.662 ;
      RECT 4.005 -28.145 4.145 -27.975 ;
      RECT 4.005 -27.248 4.095 -26.241 ;
      RECT 4.005 -26.935 4.145 -26.765 ;
      RECT 4.005 -25.439 4.095 -24.432 ;
      RECT 4.005 -24.915 4.145 -24.745 ;
      RECT 4.005 -24.018 4.095 -23.011 ;
      RECT 4.005 -23.705 4.145 -23.535 ;
      RECT 4.005 -22.209 4.095 -21.202 ;
      RECT 4.005 -21.685 4.145 -21.515 ;
      RECT 4.005 -20.788 4.095 -19.781 ;
      RECT 4.005 -20.475 4.145 -20.305 ;
      RECT 4.005 -18.979 4.095 -17.972 ;
      RECT 4.005 -18.455 4.145 -18.285 ;
      RECT 4.005 -17.558 4.095 -16.551 ;
      RECT 4.005 -17.245 4.145 -17.075 ;
      RECT 4.005 -15.749 4.095 -14.742 ;
      RECT 4.005 -15.225 4.145 -15.055 ;
      RECT 4.005 -14.328 4.095 -13.321 ;
      RECT 4.005 -14.015 4.145 -13.845 ;
      RECT 4.005 -12.519 4.095 -11.512 ;
      RECT 4.005 -11.995 4.145 -11.825 ;
      RECT 4.005 -11.098 4.095 -10.091 ;
      RECT 4.005 -10.785 4.145 -10.615 ;
      RECT 4.005 -9.289 4.095 -8.282 ;
      RECT 4.005 -8.765 4.145 -8.595 ;
      RECT 4.005 -7.868 4.095 -6.861 ;
      RECT 4.005 -7.555 4.145 -7.385 ;
      RECT 4.005 -6.059 4.095 -5.052 ;
      RECT 4.005 -5.535 4.145 -5.365 ;
      RECT 4.005 -4.638 4.095 -3.631 ;
      RECT 4.005 -4.325 4.145 -4.155 ;
      RECT 4.005 -2.829 4.095 -1.822 ;
      RECT 4.005 -2.305 4.145 -2.135 ;
      RECT 4.005 -1.408 4.095 -0.401 ;
      RECT 4.005 -1.095 4.145 -0.925 ;
      RECT 4.005 0.401 4.095 1.408 ;
      RECT 4.005 0.925 4.145 1.095 ;
      RECT 3.335 -59.815 3.505 -59.705 ;
      RECT 0.185 -59.815 3.505 -59.715 ;
      RECT 3.205 -49.858 3.295 -48.85 ;
      RECT 3.155 -49.255 3.295 -49.085 ;
      RECT 3.205 -48.05 3.295 -47.042 ;
      RECT 3.155 -47.815 3.295 -47.645 ;
      RECT 3.205 -46.628 3.295 -45.62 ;
      RECT 3.155 -46.025 3.295 -45.855 ;
      RECT 3.205 -44.82 3.295 -43.812 ;
      RECT 3.155 -44.585 3.295 -44.415 ;
      RECT 3.205 -43.398 3.295 -42.39 ;
      RECT 3.155 -42.795 3.295 -42.625 ;
      RECT 3.205 -41.59 3.295 -40.582 ;
      RECT 3.155 -41.355 3.295 -41.185 ;
      RECT 3.205 -40.168 3.295 -39.16 ;
      RECT 3.155 -39.565 3.295 -39.395 ;
      RECT 3.205 -38.36 3.295 -37.352 ;
      RECT 3.155 -38.125 3.295 -37.955 ;
      RECT 3.205 -36.938 3.295 -35.93 ;
      RECT 3.155 -36.335 3.295 -36.165 ;
      RECT 3.205 -35.13 3.295 -34.122 ;
      RECT 3.155 -34.895 3.295 -34.725 ;
      RECT 3.205 -33.708 3.295 -32.7 ;
      RECT 3.155 -33.105 3.295 -32.935 ;
      RECT 3.205 -31.9 3.295 -30.892 ;
      RECT 3.155 -31.665 3.295 -31.495 ;
      RECT 3.205 -30.478 3.295 -29.47 ;
      RECT 3.155 -29.875 3.295 -29.705 ;
      RECT 3.205 -28.67 3.295 -27.662 ;
      RECT 3.155 -28.435 3.295 -28.265 ;
      RECT 3.205 -27.248 3.295 -26.24 ;
      RECT 3.155 -26.645 3.295 -26.475 ;
      RECT 3.205 -25.44 3.295 -24.432 ;
      RECT 3.155 -25.205 3.295 -25.035 ;
      RECT 3.205 -24.018 3.295 -23.01 ;
      RECT 3.155 -23.415 3.295 -23.245 ;
      RECT 3.205 -22.21 3.295 -21.202 ;
      RECT 3.155 -21.975 3.295 -21.805 ;
      RECT 3.205 -20.788 3.295 -19.78 ;
      RECT 3.155 -20.185 3.295 -20.015 ;
      RECT 3.205 -18.98 3.295 -17.972 ;
      RECT 3.155 -18.745 3.295 -18.575 ;
      RECT 3.205 -17.558 3.295 -16.55 ;
      RECT 3.155 -16.955 3.295 -16.785 ;
      RECT 3.205 -15.75 3.295 -14.742 ;
      RECT 3.155 -15.515 3.295 -15.345 ;
      RECT 3.205 -14.328 3.295 -13.32 ;
      RECT 3.155 -13.725 3.295 -13.555 ;
      RECT 3.205 -12.52 3.295 -11.512 ;
      RECT 3.155 -12.285 3.295 -12.115 ;
      RECT 3.205 -11.098 3.295 -10.09 ;
      RECT 3.155 -10.495 3.295 -10.325 ;
      RECT 3.205 -9.29 3.295 -8.282 ;
      RECT 3.155 -9.055 3.295 -8.885 ;
      RECT 3.205 -7.868 3.295 -6.86 ;
      RECT 3.155 -7.265 3.295 -7.095 ;
      RECT 3.205 -6.06 3.295 -5.052 ;
      RECT 3.155 -5.825 3.295 -5.655 ;
      RECT 3.205 -4.638 3.295 -3.63 ;
      RECT 3.155 -4.035 3.295 -3.865 ;
      RECT 3.205 -2.83 3.295 -1.822 ;
      RECT 3.155 -2.595 3.295 -2.425 ;
      RECT 3.205 -1.408 3.295 -0.4 ;
      RECT 3.155 -0.805 3.295 -0.635 ;
      RECT 3.205 0.4 3.295 1.408 ;
      RECT 3.155 0.635 3.295 0.805 ;
      RECT 2.805 -49.858 2.895 -48.851 ;
      RECT 2.805 -49.545 2.945 -49.375 ;
      RECT 2.805 -48.049 2.895 -47.042 ;
      RECT 2.805 -47.525 2.945 -47.355 ;
      RECT 2.805 -46.628 2.895 -45.621 ;
      RECT 2.805 -46.315 2.945 -46.145 ;
      RECT 2.805 -44.819 2.895 -43.812 ;
      RECT 2.805 -44.295 2.945 -44.125 ;
      RECT 2.805 -43.398 2.895 -42.391 ;
      RECT 2.805 -43.085 2.945 -42.915 ;
      RECT 2.805 -41.589 2.895 -40.582 ;
      RECT 2.805 -41.065 2.945 -40.895 ;
      RECT 2.805 -40.168 2.895 -39.161 ;
      RECT 2.805 -39.855 2.945 -39.685 ;
      RECT 2.805 -38.359 2.895 -37.352 ;
      RECT 2.805 -37.835 2.945 -37.665 ;
      RECT 2.805 -36.938 2.895 -35.931 ;
      RECT 2.805 -36.625 2.945 -36.455 ;
      RECT 2.805 -35.129 2.895 -34.122 ;
      RECT 2.805 -34.605 2.945 -34.435 ;
      RECT 2.805 -33.708 2.895 -32.701 ;
      RECT 2.805 -33.395 2.945 -33.225 ;
      RECT 2.805 -31.899 2.895 -30.892 ;
      RECT 2.805 -31.375 2.945 -31.205 ;
      RECT 2.805 -30.478 2.895 -29.471 ;
      RECT 2.805 -30.165 2.945 -29.995 ;
      RECT 2.805 -28.669 2.895 -27.662 ;
      RECT 2.805 -28.145 2.945 -27.975 ;
      RECT 2.805 -27.248 2.895 -26.241 ;
      RECT 2.805 -26.935 2.945 -26.765 ;
      RECT 2.805 -25.439 2.895 -24.432 ;
      RECT 2.805 -24.915 2.945 -24.745 ;
      RECT 2.805 -24.018 2.895 -23.011 ;
      RECT 2.805 -23.705 2.945 -23.535 ;
      RECT 2.805 -22.209 2.895 -21.202 ;
      RECT 2.805 -21.685 2.945 -21.515 ;
      RECT 2.805 -20.788 2.895 -19.781 ;
      RECT 2.805 -20.475 2.945 -20.305 ;
      RECT 2.805 -18.979 2.895 -17.972 ;
      RECT 2.805 -18.455 2.945 -18.285 ;
      RECT 2.805 -17.558 2.895 -16.551 ;
      RECT 2.805 -17.245 2.945 -17.075 ;
      RECT 2.805 -15.749 2.895 -14.742 ;
      RECT 2.805 -15.225 2.945 -15.055 ;
      RECT 2.805 -14.328 2.895 -13.321 ;
      RECT 2.805 -14.015 2.945 -13.845 ;
      RECT 2.805 -12.519 2.895 -11.512 ;
      RECT 2.805 -11.995 2.945 -11.825 ;
      RECT 2.805 -11.098 2.895 -10.091 ;
      RECT 2.805 -10.785 2.945 -10.615 ;
      RECT 2.805 -9.289 2.895 -8.282 ;
      RECT 2.805 -8.765 2.945 -8.595 ;
      RECT 2.805 -7.868 2.895 -6.861 ;
      RECT 2.805 -7.555 2.945 -7.385 ;
      RECT 2.805 -6.059 2.895 -5.052 ;
      RECT 2.805 -5.535 2.945 -5.365 ;
      RECT 2.805 -4.638 2.895 -3.631 ;
      RECT 2.805 -4.325 2.945 -4.155 ;
      RECT 2.805 -2.829 2.895 -1.822 ;
      RECT 2.805 -2.305 2.945 -2.135 ;
      RECT 2.805 -1.408 2.895 -0.401 ;
      RECT 2.805 -1.095 2.945 -0.925 ;
      RECT 2.805 0.401 2.895 1.408 ;
      RECT 2.805 0.925 2.945 1.095 ;
      RECT 0.955 -60.005 2.435 -59.905 ;
      RECT 0.955 -60.375 1.055 -59.905 ;
      RECT 0.76 -62.715 2.335 -62.595 ;
      RECT 2.235 -63.215 2.335 -62.595 ;
      RECT 1.64 -63.215 1.74 -62.595 ;
      RECT 0.76 -63.17 0.86 -62.595 ;
      RECT 2.005 -49.858 2.095 -48.85 ;
      RECT 1.955 -49.255 2.095 -49.085 ;
      RECT 2.005 -48.05 2.095 -47.042 ;
      RECT 1.955 -47.815 2.095 -47.645 ;
      RECT 2.005 -46.628 2.095 -45.62 ;
      RECT 1.955 -46.025 2.095 -45.855 ;
      RECT 2.005 -44.82 2.095 -43.812 ;
      RECT 1.955 -44.585 2.095 -44.415 ;
      RECT 2.005 -43.398 2.095 -42.39 ;
      RECT 1.955 -42.795 2.095 -42.625 ;
      RECT 2.005 -41.59 2.095 -40.582 ;
      RECT 1.955 -41.355 2.095 -41.185 ;
      RECT 2.005 -40.168 2.095 -39.16 ;
      RECT 1.955 -39.565 2.095 -39.395 ;
      RECT 2.005 -38.36 2.095 -37.352 ;
      RECT 1.955 -38.125 2.095 -37.955 ;
      RECT 2.005 -36.938 2.095 -35.93 ;
      RECT 1.955 -36.335 2.095 -36.165 ;
      RECT 2.005 -35.13 2.095 -34.122 ;
      RECT 1.955 -34.895 2.095 -34.725 ;
      RECT 2.005 -33.708 2.095 -32.7 ;
      RECT 1.955 -33.105 2.095 -32.935 ;
      RECT 2.005 -31.9 2.095 -30.892 ;
      RECT 1.955 -31.665 2.095 -31.495 ;
      RECT 2.005 -30.478 2.095 -29.47 ;
      RECT 1.955 -29.875 2.095 -29.705 ;
      RECT 2.005 -28.67 2.095 -27.662 ;
      RECT 1.955 -28.435 2.095 -28.265 ;
      RECT 2.005 -27.248 2.095 -26.24 ;
      RECT 1.955 -26.645 2.095 -26.475 ;
      RECT 2.005 -25.44 2.095 -24.432 ;
      RECT 1.955 -25.205 2.095 -25.035 ;
      RECT 2.005 -24.018 2.095 -23.01 ;
      RECT 1.955 -23.415 2.095 -23.245 ;
      RECT 2.005 -22.21 2.095 -21.202 ;
      RECT 1.955 -21.975 2.095 -21.805 ;
      RECT 2.005 -20.788 2.095 -19.78 ;
      RECT 1.955 -20.185 2.095 -20.015 ;
      RECT 2.005 -18.98 2.095 -17.972 ;
      RECT 1.955 -18.745 2.095 -18.575 ;
      RECT 2.005 -17.558 2.095 -16.55 ;
      RECT 1.955 -16.955 2.095 -16.785 ;
      RECT 2.005 -15.75 2.095 -14.742 ;
      RECT 1.955 -15.515 2.095 -15.345 ;
      RECT 2.005 -14.328 2.095 -13.32 ;
      RECT 1.955 -13.725 2.095 -13.555 ;
      RECT 2.005 -12.52 2.095 -11.512 ;
      RECT 1.955 -12.285 2.095 -12.115 ;
      RECT 2.005 -11.098 2.095 -10.09 ;
      RECT 1.955 -10.495 2.095 -10.325 ;
      RECT 2.005 -9.29 2.095 -8.282 ;
      RECT 1.955 -9.055 2.095 -8.885 ;
      RECT 2.005 -7.868 2.095 -6.86 ;
      RECT 1.955 -7.265 2.095 -7.095 ;
      RECT 2.005 -6.06 2.095 -5.052 ;
      RECT 1.955 -5.825 2.095 -5.655 ;
      RECT 2.005 -4.638 2.095 -3.63 ;
      RECT 1.955 -4.035 2.095 -3.865 ;
      RECT 2.005 -2.83 2.095 -1.822 ;
      RECT 1.955 -2.595 2.095 -2.425 ;
      RECT 2.005 -1.408 2.095 -0.4 ;
      RECT 1.955 -0.805 2.095 -0.635 ;
      RECT 2.005 0.4 2.095 1.408 ;
      RECT 1.955 0.635 2.095 0.805 ;
      RECT 1.88 -63.005 2.055 -62.835 ;
      RECT 1.955 -63.215 2.055 -62.835 ;
      RECT 0.995 -61.875 1.095 -61.41 ;
      RECT 1.36 -61.875 1.46 -61.42 ;
      RECT 0.995 -61.875 1.84 -61.705 ;
      RECT 1.605 -49.858 1.695 -48.851 ;
      RECT 1.605 -49.545 1.745 -49.375 ;
      RECT 1.605 -48.049 1.695 -47.042 ;
      RECT 1.605 -47.525 1.745 -47.355 ;
      RECT 1.605 -46.628 1.695 -45.621 ;
      RECT 1.605 -46.315 1.745 -46.145 ;
      RECT 1.605 -44.819 1.695 -43.812 ;
      RECT 1.605 -44.295 1.745 -44.125 ;
      RECT 1.605 -43.398 1.695 -42.391 ;
      RECT 1.605 -43.085 1.745 -42.915 ;
      RECT 1.605 -41.589 1.695 -40.582 ;
      RECT 1.605 -41.065 1.745 -40.895 ;
      RECT 1.605 -40.168 1.695 -39.161 ;
      RECT 1.605 -39.855 1.745 -39.685 ;
      RECT 1.605 -38.359 1.695 -37.352 ;
      RECT 1.605 -37.835 1.745 -37.665 ;
      RECT 1.605 -36.938 1.695 -35.931 ;
      RECT 1.605 -36.625 1.745 -36.455 ;
      RECT 1.605 -35.129 1.695 -34.122 ;
      RECT 1.605 -34.605 1.745 -34.435 ;
      RECT 1.605 -33.708 1.695 -32.701 ;
      RECT 1.605 -33.395 1.745 -33.225 ;
      RECT 1.605 -31.899 1.695 -30.892 ;
      RECT 1.605 -31.375 1.745 -31.205 ;
      RECT 1.605 -30.478 1.695 -29.471 ;
      RECT 1.605 -30.165 1.745 -29.995 ;
      RECT 1.605 -28.669 1.695 -27.662 ;
      RECT 1.605 -28.145 1.745 -27.975 ;
      RECT 1.605 -27.248 1.695 -26.241 ;
      RECT 1.605 -26.935 1.745 -26.765 ;
      RECT 1.605 -25.439 1.695 -24.432 ;
      RECT 1.605 -24.915 1.745 -24.745 ;
      RECT 1.605 -24.018 1.695 -23.011 ;
      RECT 1.605 -23.705 1.745 -23.535 ;
      RECT 1.605 -22.209 1.695 -21.202 ;
      RECT 1.605 -21.685 1.745 -21.515 ;
      RECT 1.605 -20.788 1.695 -19.781 ;
      RECT 1.605 -20.475 1.745 -20.305 ;
      RECT 1.605 -18.979 1.695 -17.972 ;
      RECT 1.605 -18.455 1.745 -18.285 ;
      RECT 1.605 -17.558 1.695 -16.551 ;
      RECT 1.605 -17.245 1.745 -17.075 ;
      RECT 1.605 -15.749 1.695 -14.742 ;
      RECT 1.605 -15.225 1.745 -15.055 ;
      RECT 1.605 -14.328 1.695 -13.321 ;
      RECT 1.605 -14.015 1.745 -13.845 ;
      RECT 1.605 -12.519 1.695 -11.512 ;
      RECT 1.605 -11.995 1.745 -11.825 ;
      RECT 1.605 -11.098 1.695 -10.091 ;
      RECT 1.605 -10.785 1.745 -10.615 ;
      RECT 1.605 -9.289 1.695 -8.282 ;
      RECT 1.605 -8.765 1.745 -8.595 ;
      RECT 1.605 -7.868 1.695 -6.861 ;
      RECT 1.605 -7.555 1.745 -7.385 ;
      RECT 1.605 -6.059 1.695 -5.052 ;
      RECT 1.605 -5.535 1.745 -5.365 ;
      RECT 1.605 -4.638 1.695 -3.631 ;
      RECT 1.605 -4.325 1.745 -4.155 ;
      RECT 1.605 -2.829 1.695 -1.822 ;
      RECT 1.605 -2.305 1.745 -2.135 ;
      RECT 1.605 -1.408 1.695 -0.401 ;
      RECT 1.605 -1.095 1.745 -0.925 ;
      RECT 1.605 0.401 1.695 1.408 ;
      RECT 1.605 0.925 1.745 1.095 ;
      RECT 1.29 -63.005 1.46 -62.835 ;
      RECT 1.36 -63.215 1.46 -62.835 ;
      RECT 0.805 -49.858 0.895 -48.85 ;
      RECT 0.755 -49.255 0.895 -49.085 ;
      RECT 0.805 -48.05 0.895 -47.042 ;
      RECT 0.755 -47.815 0.895 -47.645 ;
      RECT 0.805 -46.628 0.895 -45.62 ;
      RECT 0.755 -46.025 0.895 -45.855 ;
      RECT 0.805 -44.82 0.895 -43.812 ;
      RECT 0.755 -44.585 0.895 -44.415 ;
      RECT 0.805 -43.398 0.895 -42.39 ;
      RECT 0.755 -42.795 0.895 -42.625 ;
      RECT 0.805 -41.59 0.895 -40.582 ;
      RECT 0.755 -41.355 0.895 -41.185 ;
      RECT 0.805 -40.168 0.895 -39.16 ;
      RECT 0.755 -39.565 0.895 -39.395 ;
      RECT 0.805 -38.36 0.895 -37.352 ;
      RECT 0.755 -38.125 0.895 -37.955 ;
      RECT 0.805 -36.938 0.895 -35.93 ;
      RECT 0.755 -36.335 0.895 -36.165 ;
      RECT 0.805 -35.13 0.895 -34.122 ;
      RECT 0.755 -34.895 0.895 -34.725 ;
      RECT 0.805 -33.708 0.895 -32.7 ;
      RECT 0.755 -33.105 0.895 -32.935 ;
      RECT 0.805 -31.9 0.895 -30.892 ;
      RECT 0.755 -31.665 0.895 -31.495 ;
      RECT 0.805 -30.478 0.895 -29.47 ;
      RECT 0.755 -29.875 0.895 -29.705 ;
      RECT 0.805 -28.67 0.895 -27.662 ;
      RECT 0.755 -28.435 0.895 -28.265 ;
      RECT 0.805 -27.248 0.895 -26.24 ;
      RECT 0.755 -26.645 0.895 -26.475 ;
      RECT 0.805 -25.44 0.895 -24.432 ;
      RECT 0.755 -25.205 0.895 -25.035 ;
      RECT 0.805 -24.018 0.895 -23.01 ;
      RECT 0.755 -23.415 0.895 -23.245 ;
      RECT 0.805 -22.21 0.895 -21.202 ;
      RECT 0.755 -21.975 0.895 -21.805 ;
      RECT 0.805 -20.788 0.895 -19.78 ;
      RECT 0.755 -20.185 0.895 -20.015 ;
      RECT 0.805 -18.98 0.895 -17.972 ;
      RECT 0.755 -18.745 0.895 -18.575 ;
      RECT 0.805 -17.558 0.895 -16.55 ;
      RECT 0.755 -16.955 0.895 -16.785 ;
      RECT 0.805 -15.75 0.895 -14.742 ;
      RECT 0.755 -15.515 0.895 -15.345 ;
      RECT 0.805 -14.328 0.895 -13.32 ;
      RECT 0.755 -13.725 0.895 -13.555 ;
      RECT 0.805 -12.52 0.895 -11.512 ;
      RECT 0.755 -12.285 0.895 -12.115 ;
      RECT 0.805 -11.098 0.895 -10.09 ;
      RECT 0.755 -10.495 0.895 -10.325 ;
      RECT 0.805 -9.29 0.895 -8.282 ;
      RECT 0.755 -9.055 0.895 -8.885 ;
      RECT 0.805 -7.868 0.895 -6.86 ;
      RECT 0.755 -7.265 0.895 -7.095 ;
      RECT 0.805 -6.06 0.895 -5.052 ;
      RECT 0.755 -5.825 0.895 -5.655 ;
      RECT 0.805 -4.638 0.895 -3.63 ;
      RECT 0.755 -4.035 0.895 -3.865 ;
      RECT 0.805 -2.83 0.895 -1.822 ;
      RECT 0.755 -2.595 0.895 -2.425 ;
      RECT 0.805 -1.408 0.895 -0.4 ;
      RECT 0.755 -0.805 0.895 -0.635 ;
      RECT 0.805 0.4 0.895 1.408 ;
      RECT 0.755 0.635 0.895 0.805 ;
      RECT 0.405 -49.858 0.495 -48.851 ;
      RECT 0.405 -49.545 0.545 -49.375 ;
      RECT 0.405 -48.049 0.495 -47.042 ;
      RECT 0.405 -47.525 0.545 -47.355 ;
      RECT 0.405 -46.628 0.495 -45.621 ;
      RECT 0.405 -46.315 0.545 -46.145 ;
      RECT 0.405 -44.819 0.495 -43.812 ;
      RECT 0.405 -44.295 0.545 -44.125 ;
      RECT 0.405 -43.398 0.495 -42.391 ;
      RECT 0.405 -43.085 0.545 -42.915 ;
      RECT 0.405 -41.589 0.495 -40.582 ;
      RECT 0.405 -41.065 0.545 -40.895 ;
      RECT 0.405 -40.168 0.495 -39.161 ;
      RECT 0.405 -39.855 0.545 -39.685 ;
      RECT 0.405 -38.359 0.495 -37.352 ;
      RECT 0.405 -37.835 0.545 -37.665 ;
      RECT 0.405 -36.938 0.495 -35.931 ;
      RECT 0.405 -36.625 0.545 -36.455 ;
      RECT 0.405 -35.129 0.495 -34.122 ;
      RECT 0.405 -34.605 0.545 -34.435 ;
      RECT 0.405 -33.708 0.495 -32.701 ;
      RECT 0.405 -33.395 0.545 -33.225 ;
      RECT 0.405 -31.899 0.495 -30.892 ;
      RECT 0.405 -31.375 0.545 -31.205 ;
      RECT 0.405 -30.478 0.495 -29.471 ;
      RECT 0.405 -30.165 0.545 -29.995 ;
      RECT 0.405 -28.669 0.495 -27.662 ;
      RECT 0.405 -28.145 0.545 -27.975 ;
      RECT 0.405 -27.248 0.495 -26.241 ;
      RECT 0.405 -26.935 0.545 -26.765 ;
      RECT 0.405 -25.439 0.495 -24.432 ;
      RECT 0.405 -24.915 0.545 -24.745 ;
      RECT 0.405 -24.018 0.495 -23.011 ;
      RECT 0.405 -23.705 0.545 -23.535 ;
      RECT 0.405 -22.209 0.495 -21.202 ;
      RECT 0.405 -21.685 0.545 -21.515 ;
      RECT 0.405 -20.788 0.495 -19.781 ;
      RECT 0.405 -20.475 0.545 -20.305 ;
      RECT 0.405 -18.979 0.495 -17.972 ;
      RECT 0.405 -18.455 0.545 -18.285 ;
      RECT 0.405 -17.558 0.495 -16.551 ;
      RECT 0.405 -17.245 0.545 -17.075 ;
      RECT 0.405 -15.749 0.495 -14.742 ;
      RECT 0.405 -15.225 0.545 -15.055 ;
      RECT 0.405 -14.328 0.495 -13.321 ;
      RECT 0.405 -14.015 0.545 -13.845 ;
      RECT 0.405 -12.519 0.495 -11.512 ;
      RECT 0.405 -11.995 0.545 -11.825 ;
      RECT 0.405 -11.098 0.495 -10.091 ;
      RECT 0.405 -10.785 0.545 -10.615 ;
      RECT 0.405 -9.289 0.495 -8.282 ;
      RECT 0.405 -8.765 0.545 -8.595 ;
      RECT 0.405 -7.868 0.495 -6.861 ;
      RECT 0.405 -7.555 0.545 -7.385 ;
      RECT 0.405 -6.059 0.495 -5.052 ;
      RECT 0.405 -5.535 0.545 -5.365 ;
      RECT 0.405 -4.638 0.495 -3.631 ;
      RECT 0.405 -4.325 0.545 -4.155 ;
      RECT 0.405 -2.829 0.495 -1.822 ;
      RECT 0.405 -2.305 0.545 -2.135 ;
      RECT 0.405 -1.408 0.495 -0.401 ;
      RECT 0.405 -1.095 0.545 -0.925 ;
      RECT 0.405 0.401 0.495 1.408 ;
      RECT 0.405 0.925 0.545 1.095 ;
      RECT -5.605 4.135 -5.435 4.76 ;
      RECT -6.165 4.135 -6.065 4.76 ;
      RECT -6.165 4.135 -0.245 4.235 ;
      RECT -6.165 2.91 -5.435 3.03 ;
      RECT -5.605 2.22 -5.435 3.03 ;
      RECT -6.165 2.22 -6.065 3.03 ;
      RECT -6.485 -51.435 -6.385 -50.615 ;
      RECT -7.005 -51.435 -6.905 -50.615 ;
      RECT -7.005 -51.435 -5.96 -51.335 ;
      RECT -7.005 -48.795 -5.96 -48.695 ;
      RECT -6.485 -49.515 -6.385 -48.695 ;
      RECT -7.005 -49.515 -6.905 -48.695 ;
      RECT -6.485 -38.515 -6.385 -37.695 ;
      RECT -7.005 -38.515 -6.905 -37.695 ;
      RECT -7.005 -38.515 -5.96 -38.415 ;
      RECT -7.005 -35.875 -5.96 -35.775 ;
      RECT -6.485 -36.595 -6.385 -35.775 ;
      RECT -7.005 -36.595 -6.905 -35.775 ;
      RECT -6.485 -25.595 -6.385 -24.775 ;
      RECT -7.005 -25.595 -6.905 -24.775 ;
      RECT -7.005 -25.595 -5.96 -25.495 ;
      RECT -7.005 -22.955 -5.96 -22.855 ;
      RECT -6.485 -23.675 -6.385 -22.855 ;
      RECT -7.005 -23.675 -6.905 -22.855 ;
      RECT -6.485 -12.675 -6.385 -11.855 ;
      RECT -7.005 -12.675 -6.905 -11.855 ;
      RECT -7.005 -12.675 -5.96 -12.575 ;
      RECT -7.005 -10.035 -5.96 -9.935 ;
      RECT -6.485 -10.755 -6.385 -9.935 ;
      RECT -7.005 -10.755 -6.905 -9.935 ;
      RECT -6.485 0.245 -6.385 1.065 ;
      RECT -7.005 0.245 -6.905 1.065 ;
      RECT -7.005 0.245 -5.96 0.345 ;
      RECT -7.785 -51.435 -7.685 -50.615 ;
      RECT -8.305 -51.435 -8.205 -50.615 ;
      RECT -8.305 -51.435 -7.26 -51.335 ;
      RECT -8.305 -48.795 -7.26 -48.695 ;
      RECT -7.785 -49.515 -7.685 -48.695 ;
      RECT -8.305 -49.515 -8.205 -48.695 ;
      RECT -7.785 -38.515 -7.685 -37.695 ;
      RECT -8.305 -38.515 -8.205 -37.695 ;
      RECT -8.305 -38.515 -7.26 -38.415 ;
      RECT -8.305 -35.875 -7.26 -35.775 ;
      RECT -7.785 -36.595 -7.685 -35.775 ;
      RECT -8.305 -36.595 -8.205 -35.775 ;
      RECT -7.785 -25.595 -7.685 -24.775 ;
      RECT -8.305 -25.595 -8.205 -24.775 ;
      RECT -8.305 -25.595 -7.26 -25.495 ;
      RECT -8.305 -22.955 -7.26 -22.855 ;
      RECT -7.785 -23.675 -7.685 -22.855 ;
      RECT -8.305 -23.675 -8.205 -22.855 ;
      RECT -7.785 -12.675 -7.685 -11.855 ;
      RECT -8.305 -12.675 -8.205 -11.855 ;
      RECT -8.305 -12.675 -7.26 -12.575 ;
      RECT -8.305 -10.035 -7.26 -9.935 ;
      RECT -7.785 -10.755 -7.685 -9.935 ;
      RECT -8.305 -10.755 -8.205 -9.935 ;
      RECT -7.785 0.245 -7.685 1.065 ;
      RECT -8.305 0.245 -8.205 1.065 ;
      RECT -8.305 0.245 -7.26 0.345 ;
      RECT -9.085 -51.435 -8.985 -50.615 ;
      RECT -9.605 -51.435 -9.505 -50.615 ;
      RECT -9.605 -51.435 -8.56 -51.335 ;
      RECT -9.605 -48.795 -8.56 -48.695 ;
      RECT -9.085 -49.515 -8.985 -48.695 ;
      RECT -9.605 -49.515 -9.505 -48.695 ;
      RECT -9.085 -38.515 -8.985 -37.695 ;
      RECT -9.605 -38.515 -9.505 -37.695 ;
      RECT -9.605 -38.515 -8.56 -38.415 ;
      RECT -9.605 -35.875 -8.56 -35.775 ;
      RECT -9.085 -36.595 -8.985 -35.775 ;
      RECT -9.605 -36.595 -9.505 -35.775 ;
      RECT -9.085 -25.595 -8.985 -24.775 ;
      RECT -9.605 -25.595 -9.505 -24.775 ;
      RECT -9.605 -25.595 -8.56 -25.495 ;
      RECT -9.605 -22.955 -8.56 -22.855 ;
      RECT -9.085 -23.675 -8.985 -22.855 ;
      RECT -9.605 -23.675 -9.505 -22.855 ;
      RECT -9.085 -12.675 -8.985 -11.855 ;
      RECT -9.605 -12.675 -9.505 -11.855 ;
      RECT -9.605 -12.675 -8.56 -12.575 ;
      RECT -9.605 -10.035 -8.56 -9.935 ;
      RECT -9.085 -10.755 -8.985 -9.935 ;
      RECT -9.605 -10.755 -9.505 -9.935 ;
      RECT -9.085 0.245 -8.985 1.065 ;
      RECT -9.605 0.245 -9.505 1.065 ;
      RECT -9.605 0.245 -8.56 0.345 ;
      RECT -10.385 -51.435 -10.285 -50.615 ;
      RECT -10.905 -51.435 -10.805 -50.615 ;
      RECT -10.905 -51.435 -9.86 -51.335 ;
      RECT -10.905 -48.795 -9.86 -48.695 ;
      RECT -10.385 -49.515 -10.285 -48.695 ;
      RECT -10.905 -49.515 -10.805 -48.695 ;
      RECT -10.385 -38.515 -10.285 -37.695 ;
      RECT -10.905 -38.515 -10.805 -37.695 ;
      RECT -10.905 -38.515 -9.86 -38.415 ;
      RECT -10.905 -35.875 -9.86 -35.775 ;
      RECT -10.385 -36.595 -10.285 -35.775 ;
      RECT -10.905 -36.595 -10.805 -35.775 ;
      RECT -10.385 -25.595 -10.285 -24.775 ;
      RECT -10.905 -25.595 -10.805 -24.775 ;
      RECT -10.905 -25.595 -9.86 -25.495 ;
      RECT -10.905 -22.955 -9.86 -22.855 ;
      RECT -10.385 -23.675 -10.285 -22.855 ;
      RECT -10.905 -23.675 -10.805 -22.855 ;
      RECT -10.385 -12.675 -10.285 -11.855 ;
      RECT -10.905 -12.675 -10.805 -11.855 ;
      RECT -10.905 -12.675 -9.86 -12.575 ;
      RECT -10.905 -10.035 -9.86 -9.935 ;
      RECT -10.385 -10.755 -10.285 -9.935 ;
      RECT -10.905 -10.755 -10.805 -9.935 ;
      RECT -10.385 0.245 -10.285 1.065 ;
      RECT -10.905 0.245 -10.805 1.065 ;
      RECT -10.905 0.245 -9.86 0.345 ;
      RECT -12.205 -48.795 -11.16 -48.695 ;
      RECT -11.685 -49.515 -11.585 -48.695 ;
      RECT -12.205 -49.515 -12.105 -48.695 ;
      RECT -11.685 -38.515 -11.585 -37.695 ;
      RECT -12.205 -38.515 -12.105 -37.695 ;
      RECT -12.205 -38.515 -11.16 -38.415 ;
      RECT -12.205 -35.875 -11.16 -35.775 ;
      RECT -11.685 -36.595 -11.585 -35.775 ;
      RECT -12.205 -36.595 -12.105 -35.775 ;
      RECT -11.685 -25.595 -11.585 -24.775 ;
      RECT -12.205 -25.595 -12.105 -24.775 ;
      RECT -12.205 -25.595 -11.16 -25.495 ;
      RECT -12.205 -22.955 -11.16 -22.855 ;
      RECT -11.685 -23.675 -11.585 -22.855 ;
      RECT -12.205 -23.675 -12.105 -22.855 ;
      RECT -11.685 -12.675 -11.585 -11.855 ;
      RECT -12.205 -12.675 -12.105 -11.855 ;
      RECT -12.205 -12.675 -11.16 -12.575 ;
      RECT -12.205 -10.035 -11.16 -9.935 ;
      RECT -11.685 -10.755 -11.585 -9.935 ;
      RECT -12.205 -10.755 -12.105 -9.935 ;
      RECT -11.685 0.245 -11.585 1.065 ;
      RECT -12.205 0.245 -12.105 1.065 ;
      RECT -12.205 0.245 -11.16 0.345 ;
      RECT -13.505 -48.795 -12.46 -48.695 ;
      RECT -12.985 -49.515 -12.885 -48.695 ;
      RECT -13.505 -49.515 -13.405 -48.695 ;
      RECT -12.985 -38.515 -12.885 -37.695 ;
      RECT -13.505 -38.515 -13.405 -37.695 ;
      RECT -13.505 -38.515 -12.46 -38.415 ;
      RECT -13.505 -35.875 -12.46 -35.775 ;
      RECT -12.985 -36.595 -12.885 -35.775 ;
      RECT -13.505 -36.595 -13.405 -35.775 ;
      RECT -12.985 -25.595 -12.885 -24.775 ;
      RECT -13.505 -25.595 -13.405 -24.775 ;
      RECT -13.505 -25.595 -12.46 -25.495 ;
      RECT -13.505 -22.955 -12.46 -22.855 ;
      RECT -12.985 -23.675 -12.885 -22.855 ;
      RECT -13.505 -23.675 -13.405 -22.855 ;
      RECT -12.985 -12.675 -12.885 -11.855 ;
      RECT -13.505 -12.675 -13.405 -11.855 ;
      RECT -13.505 -12.675 -12.46 -12.575 ;
      RECT -13.505 -10.035 -12.46 -9.935 ;
      RECT -12.985 -10.755 -12.885 -9.935 ;
      RECT -13.505 -10.755 -13.405 -9.935 ;
      RECT -12.985 0.245 -12.885 1.065 ;
      RECT -13.505 0.245 -13.405 1.065 ;
      RECT -13.505 0.245 -12.46 0.345 ;
      RECT -14.805 -48.795 -13.76 -48.695 ;
      RECT -14.285 -49.515 -14.185 -48.695 ;
      RECT -14.805 -49.515 -14.705 -48.695 ;
      RECT -14.285 -38.515 -14.185 -37.695 ;
      RECT -14.805 -38.515 -14.705 -37.695 ;
      RECT -14.805 -38.515 -13.76 -38.415 ;
      RECT -14.805 -35.875 -13.76 -35.775 ;
      RECT -14.285 -36.595 -14.185 -35.775 ;
      RECT -14.805 -36.595 -14.705 -35.775 ;
      RECT -14.285 -25.595 -14.185 -24.775 ;
      RECT -14.805 -25.595 -14.705 -24.775 ;
      RECT -14.805 -25.595 -13.76 -25.495 ;
      RECT -14.805 -22.955 -13.76 -22.855 ;
      RECT -14.285 -23.675 -14.185 -22.855 ;
      RECT -14.805 -23.675 -14.705 -22.855 ;
      RECT -14.285 -12.675 -14.185 -11.855 ;
      RECT -14.805 -12.675 -14.705 -11.855 ;
      RECT -14.805 -12.675 -13.76 -12.575 ;
      RECT -14.805 -10.035 -13.76 -9.935 ;
      RECT -14.285 -10.755 -14.185 -9.935 ;
      RECT -14.805 -10.755 -14.705 -9.935 ;
      RECT -14.285 0.245 -14.185 1.065 ;
      RECT -14.805 0.245 -14.705 1.065 ;
      RECT -14.805 0.245 -13.76 0.345 ;
      RECT -16.105 -48.795 -15.06 -48.695 ;
      RECT -15.585 -49.515 -15.485 -48.695 ;
      RECT -16.105 -49.515 -16.005 -48.695 ;
      RECT -15.585 -38.515 -15.485 -37.695 ;
      RECT -16.105 -38.515 -16.005 -37.695 ;
      RECT -16.105 -38.515 -15.06 -38.415 ;
      RECT -16.105 -35.875 -15.06 -35.775 ;
      RECT -15.585 -36.595 -15.485 -35.775 ;
      RECT -16.105 -36.595 -16.005 -35.775 ;
      RECT -15.585 -25.595 -15.485 -24.775 ;
      RECT -16.105 -25.595 -16.005 -24.775 ;
      RECT -16.105 -25.595 -15.06 -25.495 ;
      RECT -16.105 -22.955 -15.06 -22.855 ;
      RECT -15.585 -23.675 -15.485 -22.855 ;
      RECT -16.105 -23.675 -16.005 -22.855 ;
      RECT -15.585 -12.675 -15.485 -11.855 ;
      RECT -16.105 -12.675 -16.005 -11.855 ;
      RECT -16.105 -12.675 -15.06 -12.575 ;
      RECT -16.105 -10.035 -15.06 -9.935 ;
      RECT -15.585 -10.755 -15.485 -9.935 ;
      RECT -16.105 -10.755 -16.005 -9.935 ;
      RECT -15.585 0.245 -15.485 1.065 ;
      RECT -16.105 0.245 -16.005 1.065 ;
      RECT -16.105 0.245 -15.06 0.345 ;
      RECT -17.405 -48.795 -16.36 -48.695 ;
      RECT -16.885 -49.515 -16.785 -48.695 ;
      RECT -17.405 -49.515 -17.305 -48.695 ;
      RECT -16.885 -38.515 -16.785 -37.695 ;
      RECT -17.405 -38.515 -17.305 -37.695 ;
      RECT -17.405 -38.515 -16.36 -38.415 ;
      RECT -17.405 -35.875 -16.36 -35.775 ;
      RECT -16.885 -36.595 -16.785 -35.775 ;
      RECT -17.405 -36.595 -17.305 -35.775 ;
      RECT -16.885 -25.595 -16.785 -24.775 ;
      RECT -17.405 -25.595 -17.305 -24.775 ;
      RECT -17.405 -25.595 -16.36 -25.495 ;
      RECT -17.405 -22.955 -16.36 -22.855 ;
      RECT -16.885 -23.675 -16.785 -22.855 ;
      RECT -17.405 -23.675 -17.305 -22.855 ;
      RECT -16.885 -12.675 -16.785 -11.855 ;
      RECT -17.405 -12.675 -17.305 -11.855 ;
      RECT -17.405 -12.675 -16.36 -12.575 ;
      RECT -17.405 -10.035 -16.36 -9.935 ;
      RECT -16.885 -10.755 -16.785 -9.935 ;
      RECT -17.405 -10.755 -17.305 -9.935 ;
      RECT -16.885 0.245 -16.785 1.065 ;
      RECT -17.405 0.245 -17.305 1.065 ;
      RECT -17.405 0.245 -16.36 0.345 ;
      RECT -18.705 -48.795 -17.66 -48.695 ;
      RECT -18.185 -49.515 -18.085 -48.695 ;
      RECT -18.705 -49.515 -18.605 -48.695 ;
      RECT -18.185 -38.515 -18.085 -37.695 ;
      RECT -18.705 -38.515 -18.605 -37.695 ;
      RECT -18.705 -38.515 -17.66 -38.415 ;
      RECT -18.705 -35.875 -17.66 -35.775 ;
      RECT -18.185 -36.595 -18.085 -35.775 ;
      RECT -18.705 -36.595 -18.605 -35.775 ;
      RECT -18.185 -25.595 -18.085 -24.775 ;
      RECT -18.705 -25.595 -18.605 -24.775 ;
      RECT -18.705 -25.595 -17.66 -25.495 ;
      RECT -18.705 -22.955 -17.66 -22.855 ;
      RECT -18.185 -23.675 -18.085 -22.855 ;
      RECT -18.705 -23.675 -18.605 -22.855 ;
      RECT -18.185 -12.675 -18.085 -11.855 ;
      RECT -18.705 -12.675 -18.605 -11.855 ;
      RECT -18.705 -12.675 -17.66 -12.575 ;
      RECT -18.705 -10.035 -17.66 -9.935 ;
      RECT -18.185 -10.755 -18.085 -9.935 ;
      RECT -18.705 -10.755 -18.605 -9.935 ;
      RECT -18.185 0.245 -18.085 1.065 ;
      RECT -18.705 0.245 -18.605 1.065 ;
      RECT -18.705 0.245 -17.66 0.345 ;
      RECT -20.005 -48.795 -18.96 -48.695 ;
      RECT -19.485 -49.515 -19.385 -48.695 ;
      RECT -20.005 -49.515 -19.905 -48.695 ;
      RECT -19.485 -38.515 -19.385 -37.695 ;
      RECT -20.005 -38.515 -19.905 -37.695 ;
      RECT -20.005 -38.515 -18.96 -38.415 ;
      RECT -20.005 -35.875 -18.96 -35.775 ;
      RECT -19.485 -36.595 -19.385 -35.775 ;
      RECT -20.005 -36.595 -19.905 -35.775 ;
      RECT -19.485 -25.595 -19.385 -24.775 ;
      RECT -20.005 -25.595 -19.905 -24.775 ;
      RECT -20.005 -25.595 -18.96 -25.495 ;
      RECT -20.005 -22.955 -18.96 -22.855 ;
      RECT -19.485 -23.675 -19.385 -22.855 ;
      RECT -20.005 -23.675 -19.905 -22.855 ;
      RECT -19.485 -12.675 -19.385 -11.855 ;
      RECT -20.005 -12.675 -19.905 -11.855 ;
      RECT -20.005 -12.675 -18.96 -12.575 ;
      RECT -20.005 -10.035 -18.96 -9.935 ;
      RECT -19.485 -10.755 -19.385 -9.935 ;
      RECT -20.005 -10.755 -19.905 -9.935 ;
      RECT -19.485 0.245 -19.385 1.065 ;
      RECT -20.005 0.245 -19.905 1.065 ;
      RECT -20.005 0.245 -18.96 0.345 ;
      RECT -21.305 -48.795 -20.26 -48.695 ;
      RECT -20.785 -49.515 -20.685 -48.695 ;
      RECT -21.305 -49.515 -21.205 -48.695 ;
      RECT -20.785 -38.515 -20.685 -37.695 ;
      RECT -21.305 -38.515 -21.205 -37.695 ;
      RECT -21.305 -38.515 -20.26 -38.415 ;
      RECT -21.305 -35.875 -20.26 -35.775 ;
      RECT -20.785 -36.595 -20.685 -35.775 ;
      RECT -21.305 -36.595 -21.205 -35.775 ;
      RECT -20.785 -25.595 -20.685 -24.775 ;
      RECT -21.305 -25.595 -21.205 -24.775 ;
      RECT -21.305 -25.595 -20.26 -25.495 ;
      RECT -21.305 -22.955 -20.26 -22.855 ;
      RECT -20.785 -23.675 -20.685 -22.855 ;
      RECT -21.305 -23.675 -21.205 -22.855 ;
      RECT -20.785 -12.675 -20.685 -11.855 ;
      RECT -21.305 -12.675 -21.205 -11.855 ;
      RECT -21.305 -12.675 -20.26 -12.575 ;
      RECT -21.305 -10.035 -20.26 -9.935 ;
      RECT -20.785 -10.755 -20.685 -9.935 ;
      RECT -21.305 -10.755 -21.205 -9.935 ;
      RECT -20.785 0.245 -20.685 1.065 ;
      RECT -21.305 0.245 -21.205 1.065 ;
      RECT -21.305 0.245 -20.26 0.345 ;
      RECT -22.605 -48.795 -21.56 -48.695 ;
      RECT -22.085 -49.515 -21.985 -48.695 ;
      RECT -22.605 -49.515 -22.505 -48.695 ;
      RECT -22.085 -38.515 -21.985 -37.695 ;
      RECT -22.605 -38.515 -22.505 -37.695 ;
      RECT -22.605 -38.515 -21.56 -38.415 ;
      RECT -22.605 -35.875 -21.56 -35.775 ;
      RECT -22.085 -36.595 -21.985 -35.775 ;
      RECT -22.605 -36.595 -22.505 -35.775 ;
      RECT -22.085 -25.595 -21.985 -24.775 ;
      RECT -22.605 -25.595 -22.505 -24.775 ;
      RECT -22.605 -25.595 -21.56 -25.495 ;
      RECT -22.605 -22.955 -21.56 -22.855 ;
      RECT -22.085 -23.675 -21.985 -22.855 ;
      RECT -22.605 -23.675 -22.505 -22.855 ;
      RECT -22.085 -12.675 -21.985 -11.855 ;
      RECT -22.605 -12.675 -22.505 -11.855 ;
      RECT -22.605 -12.675 -21.56 -12.575 ;
      RECT -22.605 -10.035 -21.56 -9.935 ;
      RECT -22.085 -10.755 -21.985 -9.935 ;
      RECT -22.605 -10.755 -22.505 -9.935 ;
      RECT -22.085 0.245 -21.985 1.065 ;
      RECT -22.605 0.245 -22.505 1.065 ;
      RECT -22.605 0.245 -21.56 0.345 ;
      RECT -23.905 -48.795 -22.86 -48.695 ;
      RECT -23.385 -49.515 -23.285 -48.695 ;
      RECT -23.905 -49.515 -23.805 -48.695 ;
      RECT -23.385 -38.515 -23.285 -37.695 ;
      RECT -23.905 -38.515 -23.805 -37.695 ;
      RECT -23.905 -38.515 -22.86 -38.415 ;
      RECT -23.905 -35.875 -22.86 -35.775 ;
      RECT -23.385 -36.595 -23.285 -35.775 ;
      RECT -23.905 -36.595 -23.805 -35.775 ;
      RECT -23.385 -25.595 -23.285 -24.775 ;
      RECT -23.905 -25.595 -23.805 -24.775 ;
      RECT -23.905 -25.595 -22.86 -25.495 ;
      RECT -23.905 -22.955 -22.86 -22.855 ;
      RECT -23.385 -23.675 -23.285 -22.855 ;
      RECT -23.905 -23.675 -23.805 -22.855 ;
      RECT -23.385 -12.675 -23.285 -11.855 ;
      RECT -23.905 -12.675 -23.805 -11.855 ;
      RECT -23.905 -12.675 -22.86 -12.575 ;
      RECT -23.905 -10.035 -22.86 -9.935 ;
      RECT -23.385 -10.755 -23.285 -9.935 ;
      RECT -23.905 -10.755 -23.805 -9.935 ;
      RECT -23.385 0.245 -23.285 1.065 ;
      RECT -23.905 0.245 -23.805 1.065 ;
      RECT -23.905 0.245 -22.86 0.345 ;
      RECT -25.205 -48.795 -24.16 -48.695 ;
      RECT -24.685 -49.515 -24.585 -48.695 ;
      RECT -25.205 -49.515 -25.105 -48.695 ;
      RECT -24.685 -38.515 -24.585 -37.695 ;
      RECT -25.205 -38.515 -25.105 -37.695 ;
      RECT -25.205 -38.515 -24.16 -38.415 ;
      RECT -25.205 -35.875 -24.16 -35.775 ;
      RECT -24.685 -36.595 -24.585 -35.775 ;
      RECT -25.205 -36.595 -25.105 -35.775 ;
      RECT -24.685 -25.595 -24.585 -24.775 ;
      RECT -25.205 -25.595 -25.105 -24.775 ;
      RECT -25.205 -25.595 -24.16 -25.495 ;
      RECT -25.205 -22.955 -24.16 -22.855 ;
      RECT -24.685 -23.675 -24.585 -22.855 ;
      RECT -25.205 -23.675 -25.105 -22.855 ;
      RECT -24.685 -12.675 -24.585 -11.855 ;
      RECT -25.205 -12.675 -25.105 -11.855 ;
      RECT -25.205 -12.675 -24.16 -12.575 ;
      RECT -25.205 -10.035 -24.16 -9.935 ;
      RECT -24.685 -10.755 -24.585 -9.935 ;
      RECT -25.205 -10.755 -25.105 -9.935 ;
      RECT -24.685 0.245 -24.585 1.065 ;
      RECT -25.205 0.245 -25.105 1.065 ;
      RECT -25.205 0.245 -24.16 0.345 ;
      RECT -26.505 -48.795 -25.46 -48.695 ;
      RECT -25.985 -49.515 -25.885 -48.695 ;
      RECT -26.505 -49.515 -26.405 -48.695 ;
      RECT -25.985 -38.515 -25.885 -37.695 ;
      RECT -26.505 -38.515 -26.405 -37.695 ;
      RECT -26.505 -38.515 -25.46 -38.415 ;
      RECT -26.505 -35.875 -25.46 -35.775 ;
      RECT -25.985 -36.595 -25.885 -35.775 ;
      RECT -26.505 -36.595 -26.405 -35.775 ;
      RECT -25.985 -25.595 -25.885 -24.775 ;
      RECT -26.505 -25.595 -26.405 -24.775 ;
      RECT -26.505 -25.595 -25.46 -25.495 ;
      RECT -26.505 -22.955 -25.46 -22.855 ;
      RECT -25.985 -23.675 -25.885 -22.855 ;
      RECT -26.505 -23.675 -26.405 -22.855 ;
      RECT -25.985 -12.675 -25.885 -11.855 ;
      RECT -26.505 -12.675 -26.405 -11.855 ;
      RECT -26.505 -12.675 -25.46 -12.575 ;
      RECT -26.505 -10.035 -25.46 -9.935 ;
      RECT -25.985 -10.755 -25.885 -9.935 ;
      RECT -26.505 -10.755 -26.405 -9.935 ;
      RECT -25.985 0.245 -25.885 1.065 ;
      RECT -26.505 0.245 -26.405 1.065 ;
      RECT -26.505 0.245 -25.46 0.345 ;
      RECT -0.425 1.935 38.945 2.035 ;
      RECT 38.275 -53.265 38.375 -52.305 ;
      RECT 37.9 -48.51 38.25 -48.39 ;
      RECT 37.9 -45.28 38.25 -45.16 ;
      RECT 37.9 -42.05 38.25 -41.93 ;
      RECT 37.9 -38.82 38.25 -38.7 ;
      RECT 37.9 -35.59 38.25 -35.47 ;
      RECT 37.9 -32.36 38.25 -32.24 ;
      RECT 37.9 -29.13 38.25 -29.01 ;
      RECT 37.9 -25.9 38.25 -25.78 ;
      RECT 37.9 -22.67 38.25 -22.55 ;
      RECT 37.9 -19.44 38.25 -19.32 ;
      RECT 37.9 -16.21 38.25 -16.09 ;
      RECT 37.9 -12.98 38.25 -12.86 ;
      RECT 37.9 -9.75 38.25 -9.63 ;
      RECT 37.9 -6.52 38.25 -6.4 ;
      RECT 37.9 -3.29 38.25 -3.17 ;
      RECT 37.9 -0.06 38.25 0.06 ;
      RECT 38.015 -53.265 38.115 -52.305 ;
      RECT 38.015 2.175 38.115 3.135 ;
      RECT 37.725 -60.575 37.825 -60.095 ;
      RECT 37.725 -59.085 37.825 -58.615 ;
      RECT 37.415 -48.51 37.765 -48.39 ;
      RECT 37.415 -45.28 37.765 -45.16 ;
      RECT 37.415 -42.05 37.765 -41.93 ;
      RECT 37.415 -38.82 37.765 -38.7 ;
      RECT 37.415 -35.59 37.765 -35.47 ;
      RECT 37.415 -32.36 37.765 -32.24 ;
      RECT 37.415 -29.13 37.765 -29.01 ;
      RECT 37.415 -25.9 37.765 -25.78 ;
      RECT 37.415 -22.67 37.765 -22.55 ;
      RECT 37.415 -19.44 37.765 -19.32 ;
      RECT 37.415 -16.21 37.765 -16.09 ;
      RECT 37.415 -12.98 37.765 -12.86 ;
      RECT 37.415 -9.75 37.765 -9.63 ;
      RECT 37.415 -6.52 37.765 -6.4 ;
      RECT 37.415 -3.29 37.765 -3.17 ;
      RECT 37.415 -0.06 37.765 0.06 ;
      RECT 37.585 -53.265 37.685 -52.305 ;
      RECT 37.585 2.175 37.685 3.135 ;
      RECT 33.685 -56.975 37.465 -56.855 ;
      RECT 37.325 -53.265 37.425 -52.305 ;
      RECT 37.135 -59.07 37.255 -58.69 ;
      RECT 37.135 -60.565 37.235 -60.095 ;
      RECT 37.075 -53.265 37.175 -52.305 ;
      RECT 36.7 -48.51 37.05 -48.39 ;
      RECT 36.7 -45.28 37.05 -45.16 ;
      RECT 36.7 -42.05 37.05 -41.93 ;
      RECT 36.7 -38.82 37.05 -38.7 ;
      RECT 36.7 -35.59 37.05 -35.47 ;
      RECT 36.7 -32.36 37.05 -32.24 ;
      RECT 36.7 -29.13 37.05 -29.01 ;
      RECT 36.7 -25.9 37.05 -25.78 ;
      RECT 36.7 -22.67 37.05 -22.55 ;
      RECT 36.7 -19.44 37.05 -19.32 ;
      RECT 36.7 -16.21 37.05 -16.09 ;
      RECT 36.7 -12.98 37.05 -12.86 ;
      RECT 36.7 -9.75 37.05 -9.63 ;
      RECT 36.7 -6.52 37.05 -6.4 ;
      RECT 36.7 -3.29 37.05 -3.17 ;
      RECT 36.7 -0.06 37.05 0.06 ;
      RECT 36.815 -53.265 36.915 -52.305 ;
      RECT 36.815 2.175 36.915 3.135 ;
      RECT 36.545 -57.915 36.68 -57.595 ;
      RECT 36.215 -48.51 36.565 -48.39 ;
      RECT 36.215 -45.28 36.565 -45.16 ;
      RECT 36.215 -42.05 36.565 -41.93 ;
      RECT 36.215 -38.82 36.565 -38.7 ;
      RECT 36.215 -35.59 36.565 -35.47 ;
      RECT 36.215 -32.36 36.565 -32.24 ;
      RECT 36.215 -29.13 36.565 -29.01 ;
      RECT 36.215 -25.9 36.565 -25.78 ;
      RECT 36.215 -22.67 36.565 -22.55 ;
      RECT 36.215 -19.44 36.565 -19.32 ;
      RECT 36.215 -16.21 36.565 -16.09 ;
      RECT 36.215 -12.98 36.565 -12.86 ;
      RECT 36.215 -9.75 36.565 -9.63 ;
      RECT 36.215 -6.52 36.565 -6.4 ;
      RECT 36.215 -3.29 36.565 -3.17 ;
      RECT 36.215 -0.06 36.565 0.06 ;
      RECT 36.385 -53.265 36.485 -52.305 ;
      RECT 36.385 2.175 36.485 3.135 ;
      RECT 36.21 -57.915 36.355 -57.595 ;
      RECT 36.125 -53.265 36.225 -52.305 ;
      RECT 35.875 -56.495 35.975 -55.535 ;
      RECT 35.5 -48.51 35.85 -48.39 ;
      RECT 35.5 -45.28 35.85 -45.16 ;
      RECT 35.5 -42.05 35.85 -41.93 ;
      RECT 35.5 -38.82 35.85 -38.7 ;
      RECT 35.5 -35.59 35.85 -35.47 ;
      RECT 35.5 -32.36 35.85 -32.24 ;
      RECT 35.5 -29.13 35.85 -29.01 ;
      RECT 35.5 -25.9 35.85 -25.78 ;
      RECT 35.5 -22.67 35.85 -22.55 ;
      RECT 35.5 -19.44 35.85 -19.32 ;
      RECT 35.5 -16.21 35.85 -16.09 ;
      RECT 35.5 -12.98 35.85 -12.86 ;
      RECT 35.5 -9.75 35.85 -9.63 ;
      RECT 35.5 -6.52 35.85 -6.4 ;
      RECT 35.5 -3.29 35.85 -3.17 ;
      RECT 35.5 -0.06 35.85 0.06 ;
      RECT 35.705 -60.575 35.805 -60.095 ;
      RECT 35.705 -59.085 35.805 -58.615 ;
      RECT 35.615 -56.495 35.715 -55.535 ;
      RECT 35.615 2.175 35.715 3.135 ;
      RECT 35.015 -48.51 35.365 -48.39 ;
      RECT 35.015 -45.28 35.365 -45.16 ;
      RECT 35.015 -42.05 35.365 -41.93 ;
      RECT 35.015 -38.82 35.365 -38.7 ;
      RECT 35.015 -35.59 35.365 -35.47 ;
      RECT 35.015 -32.36 35.365 -32.24 ;
      RECT 35.015 -29.13 35.365 -29.01 ;
      RECT 35.015 -25.9 35.365 -25.78 ;
      RECT 35.015 -22.67 35.365 -22.55 ;
      RECT 35.015 -19.44 35.365 -19.32 ;
      RECT 35.015 -16.21 35.365 -16.09 ;
      RECT 35.015 -12.98 35.365 -12.86 ;
      RECT 35.015 -9.75 35.365 -9.63 ;
      RECT 35.015 -6.52 35.365 -6.4 ;
      RECT 35.015 -3.29 35.365 -3.17 ;
      RECT 35.015 -0.06 35.365 0.06 ;
      RECT 35.185 -56.495 35.285 -55.535 ;
      RECT 35.185 2.175 35.285 3.135 ;
      RECT 35.08 -59.085 35.25 -58.705 ;
      RECT 35.115 -60.565 35.215 -60.095 ;
      RECT 34.925 -56.495 35.025 -55.535 ;
      RECT 34.675 -56.495 34.775 -55.535 ;
      RECT 34.3 -48.51 34.65 -48.39 ;
      RECT 34.3 -45.28 34.65 -45.16 ;
      RECT 34.3 -42.05 34.65 -41.93 ;
      RECT 34.3 -38.82 34.65 -38.7 ;
      RECT 34.3 -35.59 34.65 -35.47 ;
      RECT 34.3 -32.36 34.65 -32.24 ;
      RECT 34.3 -29.13 34.65 -29.01 ;
      RECT 34.3 -25.9 34.65 -25.78 ;
      RECT 34.3 -22.67 34.65 -22.55 ;
      RECT 34.3 -19.44 34.65 -19.32 ;
      RECT 34.3 -16.21 34.65 -16.09 ;
      RECT 34.3 -12.98 34.65 -12.86 ;
      RECT 34.3 -9.75 34.65 -9.63 ;
      RECT 34.3 -6.52 34.65 -6.4 ;
      RECT 34.3 -3.29 34.65 -3.17 ;
      RECT 34.3 -0.06 34.65 0.06 ;
      RECT 34.415 -56.495 34.515 -55.535 ;
      RECT 34.415 2.175 34.515 3.135 ;
      RECT 34.315 -61.875 34.415 -61.405 ;
      RECT 33.815 -48.51 34.165 -48.39 ;
      RECT 33.815 -45.28 34.165 -45.16 ;
      RECT 33.815 -42.05 34.165 -41.93 ;
      RECT 33.815 -38.82 34.165 -38.7 ;
      RECT 33.815 -35.59 34.165 -35.47 ;
      RECT 33.815 -32.36 34.165 -32.24 ;
      RECT 33.815 -29.13 34.165 -29.01 ;
      RECT 33.815 -25.9 34.165 -25.78 ;
      RECT 33.815 -22.67 34.165 -22.55 ;
      RECT 33.815 -19.44 34.165 -19.32 ;
      RECT 33.815 -16.21 34.165 -16.09 ;
      RECT 33.815 -12.98 34.165 -12.86 ;
      RECT 33.815 -9.75 34.165 -9.63 ;
      RECT 33.815 -6.52 34.165 -6.4 ;
      RECT 33.815 -3.29 34.165 -3.17 ;
      RECT 33.815 -0.06 34.165 0.06 ;
      RECT 33.95 -59.055 34.1 -58.765 ;
      RECT 33.985 -56.495 34.085 -55.535 ;
      RECT 33.985 2.175 34.085 3.135 ;
      RECT 33.965 -60.51 34.065 -59.97 ;
      RECT 33.725 -61.875 33.825 -61.405 ;
      RECT 33.725 -56.495 33.825 -55.535 ;
      RECT 33.475 -53.265 33.575 -52.305 ;
      RECT 33.1 -48.51 33.45 -48.39 ;
      RECT 33.1 -45.28 33.45 -45.16 ;
      RECT 33.1 -42.05 33.45 -41.93 ;
      RECT 33.1 -38.82 33.45 -38.7 ;
      RECT 33.1 -35.59 33.45 -35.47 ;
      RECT 33.1 -32.36 33.45 -32.24 ;
      RECT 33.1 -29.13 33.45 -29.01 ;
      RECT 33.1 -25.9 33.45 -25.78 ;
      RECT 33.1 -22.67 33.45 -22.55 ;
      RECT 33.1 -19.44 33.45 -19.32 ;
      RECT 33.1 -16.21 33.45 -16.09 ;
      RECT 33.1 -12.98 33.45 -12.86 ;
      RECT 33.1 -9.75 33.45 -9.63 ;
      RECT 33.1 -6.52 33.45 -6.4 ;
      RECT 33.1 -3.29 33.45 -3.17 ;
      RECT 33.1 -0.06 33.45 0.06 ;
      RECT 33.215 -53.265 33.315 -52.305 ;
      RECT 33.215 2.175 33.315 3.135 ;
      RECT 32.925 -60.575 33.025 -60.095 ;
      RECT 32.925 -59.085 33.025 -58.615 ;
      RECT 32.615 -48.51 32.965 -48.39 ;
      RECT 32.615 -45.28 32.965 -45.16 ;
      RECT 32.615 -42.05 32.965 -41.93 ;
      RECT 32.615 -38.82 32.965 -38.7 ;
      RECT 32.615 -35.59 32.965 -35.47 ;
      RECT 32.615 -32.36 32.965 -32.24 ;
      RECT 32.615 -29.13 32.965 -29.01 ;
      RECT 32.615 -25.9 32.965 -25.78 ;
      RECT 32.615 -22.67 32.965 -22.55 ;
      RECT 32.615 -19.44 32.965 -19.32 ;
      RECT 32.615 -16.21 32.965 -16.09 ;
      RECT 32.615 -12.98 32.965 -12.86 ;
      RECT 32.615 -9.75 32.965 -9.63 ;
      RECT 32.615 -6.52 32.965 -6.4 ;
      RECT 32.615 -3.29 32.965 -3.17 ;
      RECT 32.615 -0.06 32.965 0.06 ;
      RECT 32.785 -53.265 32.885 -52.305 ;
      RECT 32.785 2.175 32.885 3.135 ;
      RECT 28.885 -56.975 32.665 -56.855 ;
      RECT 32.525 -53.265 32.625 -52.305 ;
      RECT 32.335 -59.07 32.455 -58.69 ;
      RECT 32.335 -60.565 32.435 -60.095 ;
      RECT 32.275 -53.265 32.375 -52.305 ;
      RECT 31.9 -48.51 32.25 -48.39 ;
      RECT 31.9 -45.28 32.25 -45.16 ;
      RECT 31.9 -42.05 32.25 -41.93 ;
      RECT 31.9 -38.82 32.25 -38.7 ;
      RECT 31.9 -35.59 32.25 -35.47 ;
      RECT 31.9 -32.36 32.25 -32.24 ;
      RECT 31.9 -29.13 32.25 -29.01 ;
      RECT 31.9 -25.9 32.25 -25.78 ;
      RECT 31.9 -22.67 32.25 -22.55 ;
      RECT 31.9 -19.44 32.25 -19.32 ;
      RECT 31.9 -16.21 32.25 -16.09 ;
      RECT 31.9 -12.98 32.25 -12.86 ;
      RECT 31.9 -9.75 32.25 -9.63 ;
      RECT 31.9 -6.52 32.25 -6.4 ;
      RECT 31.9 -3.29 32.25 -3.17 ;
      RECT 31.9 -0.06 32.25 0.06 ;
      RECT 32.015 -53.265 32.115 -52.305 ;
      RECT 32.015 2.175 32.115 3.135 ;
      RECT 31.745 -57.915 31.88 -57.595 ;
      RECT 31.415 -48.51 31.765 -48.39 ;
      RECT 31.415 -45.28 31.765 -45.16 ;
      RECT 31.415 -42.05 31.765 -41.93 ;
      RECT 31.415 -38.82 31.765 -38.7 ;
      RECT 31.415 -35.59 31.765 -35.47 ;
      RECT 31.415 -32.36 31.765 -32.24 ;
      RECT 31.415 -29.13 31.765 -29.01 ;
      RECT 31.415 -25.9 31.765 -25.78 ;
      RECT 31.415 -22.67 31.765 -22.55 ;
      RECT 31.415 -19.44 31.765 -19.32 ;
      RECT 31.415 -16.21 31.765 -16.09 ;
      RECT 31.415 -12.98 31.765 -12.86 ;
      RECT 31.415 -9.75 31.765 -9.63 ;
      RECT 31.415 -6.52 31.765 -6.4 ;
      RECT 31.415 -3.29 31.765 -3.17 ;
      RECT 31.415 -0.06 31.765 0.06 ;
      RECT 31.585 -53.265 31.685 -52.305 ;
      RECT 31.585 2.175 31.685 3.135 ;
      RECT 31.41 -57.915 31.555 -57.595 ;
      RECT 31.325 -53.265 31.425 -52.305 ;
      RECT 31.075 -56.495 31.175 -55.535 ;
      RECT 30.7 -48.51 31.05 -48.39 ;
      RECT 30.7 -45.28 31.05 -45.16 ;
      RECT 30.7 -42.05 31.05 -41.93 ;
      RECT 30.7 -38.82 31.05 -38.7 ;
      RECT 30.7 -35.59 31.05 -35.47 ;
      RECT 30.7 -32.36 31.05 -32.24 ;
      RECT 30.7 -29.13 31.05 -29.01 ;
      RECT 30.7 -25.9 31.05 -25.78 ;
      RECT 30.7 -22.67 31.05 -22.55 ;
      RECT 30.7 -19.44 31.05 -19.32 ;
      RECT 30.7 -16.21 31.05 -16.09 ;
      RECT 30.7 -12.98 31.05 -12.86 ;
      RECT 30.7 -9.75 31.05 -9.63 ;
      RECT 30.7 -6.52 31.05 -6.4 ;
      RECT 30.7 -3.29 31.05 -3.17 ;
      RECT 30.7 -0.06 31.05 0.06 ;
      RECT 30.905 -60.575 31.005 -60.095 ;
      RECT 30.905 -59.085 31.005 -58.615 ;
      RECT 30.815 -56.495 30.915 -55.535 ;
      RECT 30.815 2.175 30.915 3.135 ;
      RECT 30.215 -48.51 30.565 -48.39 ;
      RECT 30.215 -45.28 30.565 -45.16 ;
      RECT 30.215 -42.05 30.565 -41.93 ;
      RECT 30.215 -38.82 30.565 -38.7 ;
      RECT 30.215 -35.59 30.565 -35.47 ;
      RECT 30.215 -32.36 30.565 -32.24 ;
      RECT 30.215 -29.13 30.565 -29.01 ;
      RECT 30.215 -25.9 30.565 -25.78 ;
      RECT 30.215 -22.67 30.565 -22.55 ;
      RECT 30.215 -19.44 30.565 -19.32 ;
      RECT 30.215 -16.21 30.565 -16.09 ;
      RECT 30.215 -12.98 30.565 -12.86 ;
      RECT 30.215 -9.75 30.565 -9.63 ;
      RECT 30.215 -6.52 30.565 -6.4 ;
      RECT 30.215 -3.29 30.565 -3.17 ;
      RECT 30.215 -0.06 30.565 0.06 ;
      RECT 30.385 -56.495 30.485 -55.535 ;
      RECT 30.385 2.175 30.485 3.135 ;
      RECT 30.28 -59.085 30.45 -58.705 ;
      RECT 30.315 -60.565 30.415 -60.095 ;
      RECT 30.125 -56.495 30.225 -55.535 ;
      RECT 29.875 -56.495 29.975 -55.535 ;
      RECT 29.5 -48.51 29.85 -48.39 ;
      RECT 29.5 -45.28 29.85 -45.16 ;
      RECT 29.5 -42.05 29.85 -41.93 ;
      RECT 29.5 -38.82 29.85 -38.7 ;
      RECT 29.5 -35.59 29.85 -35.47 ;
      RECT 29.5 -32.36 29.85 -32.24 ;
      RECT 29.5 -29.13 29.85 -29.01 ;
      RECT 29.5 -25.9 29.85 -25.78 ;
      RECT 29.5 -22.67 29.85 -22.55 ;
      RECT 29.5 -19.44 29.85 -19.32 ;
      RECT 29.5 -16.21 29.85 -16.09 ;
      RECT 29.5 -12.98 29.85 -12.86 ;
      RECT 29.5 -9.75 29.85 -9.63 ;
      RECT 29.5 -6.52 29.85 -6.4 ;
      RECT 29.5 -3.29 29.85 -3.17 ;
      RECT 29.5 -0.06 29.85 0.06 ;
      RECT 29.615 -56.495 29.715 -55.535 ;
      RECT 29.615 2.175 29.715 3.135 ;
      RECT 29.515 -61.875 29.615 -61.405 ;
      RECT 29.015 -48.51 29.365 -48.39 ;
      RECT 29.015 -45.28 29.365 -45.16 ;
      RECT 29.015 -42.05 29.365 -41.93 ;
      RECT 29.015 -38.82 29.365 -38.7 ;
      RECT 29.015 -35.59 29.365 -35.47 ;
      RECT 29.015 -32.36 29.365 -32.24 ;
      RECT 29.015 -29.13 29.365 -29.01 ;
      RECT 29.015 -25.9 29.365 -25.78 ;
      RECT 29.015 -22.67 29.365 -22.55 ;
      RECT 29.015 -19.44 29.365 -19.32 ;
      RECT 29.015 -16.21 29.365 -16.09 ;
      RECT 29.015 -12.98 29.365 -12.86 ;
      RECT 29.015 -9.75 29.365 -9.63 ;
      RECT 29.015 -6.52 29.365 -6.4 ;
      RECT 29.015 -3.29 29.365 -3.17 ;
      RECT 29.015 -0.06 29.365 0.06 ;
      RECT 29.15 -59.055 29.3 -58.765 ;
      RECT 29.185 -56.495 29.285 -55.535 ;
      RECT 29.185 2.175 29.285 3.135 ;
      RECT 29.165 -60.51 29.265 -59.97 ;
      RECT 28.925 -61.875 29.025 -61.405 ;
      RECT 28.925 -56.495 29.025 -55.535 ;
      RECT 28.675 -53.265 28.775 -52.305 ;
      RECT 28.3 -48.51 28.65 -48.39 ;
      RECT 28.3 -45.28 28.65 -45.16 ;
      RECT 28.3 -42.05 28.65 -41.93 ;
      RECT 28.3 -38.82 28.65 -38.7 ;
      RECT 28.3 -35.59 28.65 -35.47 ;
      RECT 28.3 -32.36 28.65 -32.24 ;
      RECT 28.3 -29.13 28.65 -29.01 ;
      RECT 28.3 -25.9 28.65 -25.78 ;
      RECT 28.3 -22.67 28.65 -22.55 ;
      RECT 28.3 -19.44 28.65 -19.32 ;
      RECT 28.3 -16.21 28.65 -16.09 ;
      RECT 28.3 -12.98 28.65 -12.86 ;
      RECT 28.3 -9.75 28.65 -9.63 ;
      RECT 28.3 -6.52 28.65 -6.4 ;
      RECT 28.3 -3.29 28.65 -3.17 ;
      RECT 28.3 -0.06 28.65 0.06 ;
      RECT 28.415 -53.265 28.515 -52.305 ;
      RECT 28.415 2.175 28.515 3.135 ;
      RECT 28.125 -60.575 28.225 -60.095 ;
      RECT 28.125 -59.085 28.225 -58.615 ;
      RECT 27.815 -48.51 28.165 -48.39 ;
      RECT 27.815 -45.28 28.165 -45.16 ;
      RECT 27.815 -42.05 28.165 -41.93 ;
      RECT 27.815 -38.82 28.165 -38.7 ;
      RECT 27.815 -35.59 28.165 -35.47 ;
      RECT 27.815 -32.36 28.165 -32.24 ;
      RECT 27.815 -29.13 28.165 -29.01 ;
      RECT 27.815 -25.9 28.165 -25.78 ;
      RECT 27.815 -22.67 28.165 -22.55 ;
      RECT 27.815 -19.44 28.165 -19.32 ;
      RECT 27.815 -16.21 28.165 -16.09 ;
      RECT 27.815 -12.98 28.165 -12.86 ;
      RECT 27.815 -9.75 28.165 -9.63 ;
      RECT 27.815 -6.52 28.165 -6.4 ;
      RECT 27.815 -3.29 28.165 -3.17 ;
      RECT 27.815 -0.06 28.165 0.06 ;
      RECT 27.985 -53.265 28.085 -52.305 ;
      RECT 27.985 2.175 28.085 3.135 ;
      RECT 24.085 -56.975 27.865 -56.855 ;
      RECT 27.725 -53.265 27.825 -52.305 ;
      RECT 27.535 -59.07 27.655 -58.69 ;
      RECT 27.535 -60.565 27.635 -60.095 ;
      RECT 27.475 -53.265 27.575 -52.305 ;
      RECT 27.1 -48.51 27.45 -48.39 ;
      RECT 27.1 -45.28 27.45 -45.16 ;
      RECT 27.1 -42.05 27.45 -41.93 ;
      RECT 27.1 -38.82 27.45 -38.7 ;
      RECT 27.1 -35.59 27.45 -35.47 ;
      RECT 27.1 -32.36 27.45 -32.24 ;
      RECT 27.1 -29.13 27.45 -29.01 ;
      RECT 27.1 -25.9 27.45 -25.78 ;
      RECT 27.1 -22.67 27.45 -22.55 ;
      RECT 27.1 -19.44 27.45 -19.32 ;
      RECT 27.1 -16.21 27.45 -16.09 ;
      RECT 27.1 -12.98 27.45 -12.86 ;
      RECT 27.1 -9.75 27.45 -9.63 ;
      RECT 27.1 -6.52 27.45 -6.4 ;
      RECT 27.1 -3.29 27.45 -3.17 ;
      RECT 27.1 -0.06 27.45 0.06 ;
      RECT 27.215 -53.265 27.315 -52.305 ;
      RECT 27.215 2.175 27.315 3.135 ;
      RECT 26.945 -57.915 27.08 -57.595 ;
      RECT 26.615 -48.51 26.965 -48.39 ;
      RECT 26.615 -45.28 26.965 -45.16 ;
      RECT 26.615 -42.05 26.965 -41.93 ;
      RECT 26.615 -38.82 26.965 -38.7 ;
      RECT 26.615 -35.59 26.965 -35.47 ;
      RECT 26.615 -32.36 26.965 -32.24 ;
      RECT 26.615 -29.13 26.965 -29.01 ;
      RECT 26.615 -25.9 26.965 -25.78 ;
      RECT 26.615 -22.67 26.965 -22.55 ;
      RECT 26.615 -19.44 26.965 -19.32 ;
      RECT 26.615 -16.21 26.965 -16.09 ;
      RECT 26.615 -12.98 26.965 -12.86 ;
      RECT 26.615 -9.75 26.965 -9.63 ;
      RECT 26.615 -6.52 26.965 -6.4 ;
      RECT 26.615 -3.29 26.965 -3.17 ;
      RECT 26.615 -0.06 26.965 0.06 ;
      RECT 26.785 -53.265 26.885 -52.305 ;
      RECT 26.785 2.175 26.885 3.135 ;
      RECT 26.61 -57.915 26.755 -57.595 ;
      RECT 26.525 -53.265 26.625 -52.305 ;
      RECT 26.275 -56.495 26.375 -55.535 ;
      RECT 25.9 -48.51 26.25 -48.39 ;
      RECT 25.9 -45.28 26.25 -45.16 ;
      RECT 25.9 -42.05 26.25 -41.93 ;
      RECT 25.9 -38.82 26.25 -38.7 ;
      RECT 25.9 -35.59 26.25 -35.47 ;
      RECT 25.9 -32.36 26.25 -32.24 ;
      RECT 25.9 -29.13 26.25 -29.01 ;
      RECT 25.9 -25.9 26.25 -25.78 ;
      RECT 25.9 -22.67 26.25 -22.55 ;
      RECT 25.9 -19.44 26.25 -19.32 ;
      RECT 25.9 -16.21 26.25 -16.09 ;
      RECT 25.9 -12.98 26.25 -12.86 ;
      RECT 25.9 -9.75 26.25 -9.63 ;
      RECT 25.9 -6.52 26.25 -6.4 ;
      RECT 25.9 -3.29 26.25 -3.17 ;
      RECT 25.9 -0.06 26.25 0.06 ;
      RECT 26.105 -60.575 26.205 -60.095 ;
      RECT 26.105 -59.085 26.205 -58.615 ;
      RECT 26.015 -56.495 26.115 -55.535 ;
      RECT 26.015 2.175 26.115 3.135 ;
      RECT 25.415 -48.51 25.765 -48.39 ;
      RECT 25.415 -45.28 25.765 -45.16 ;
      RECT 25.415 -42.05 25.765 -41.93 ;
      RECT 25.415 -38.82 25.765 -38.7 ;
      RECT 25.415 -35.59 25.765 -35.47 ;
      RECT 25.415 -32.36 25.765 -32.24 ;
      RECT 25.415 -29.13 25.765 -29.01 ;
      RECT 25.415 -25.9 25.765 -25.78 ;
      RECT 25.415 -22.67 25.765 -22.55 ;
      RECT 25.415 -19.44 25.765 -19.32 ;
      RECT 25.415 -16.21 25.765 -16.09 ;
      RECT 25.415 -12.98 25.765 -12.86 ;
      RECT 25.415 -9.75 25.765 -9.63 ;
      RECT 25.415 -6.52 25.765 -6.4 ;
      RECT 25.415 -3.29 25.765 -3.17 ;
      RECT 25.415 -0.06 25.765 0.06 ;
      RECT 25.585 -56.495 25.685 -55.535 ;
      RECT 25.585 2.175 25.685 3.135 ;
      RECT 25.48 -59.085 25.65 -58.705 ;
      RECT 25.515 -60.565 25.615 -60.095 ;
      RECT 25.325 -56.495 25.425 -55.535 ;
      RECT 25.075 -56.495 25.175 -55.535 ;
      RECT 24.7 -48.51 25.05 -48.39 ;
      RECT 24.7 -45.28 25.05 -45.16 ;
      RECT 24.7 -42.05 25.05 -41.93 ;
      RECT 24.7 -38.82 25.05 -38.7 ;
      RECT 24.7 -35.59 25.05 -35.47 ;
      RECT 24.7 -32.36 25.05 -32.24 ;
      RECT 24.7 -29.13 25.05 -29.01 ;
      RECT 24.7 -25.9 25.05 -25.78 ;
      RECT 24.7 -22.67 25.05 -22.55 ;
      RECT 24.7 -19.44 25.05 -19.32 ;
      RECT 24.7 -16.21 25.05 -16.09 ;
      RECT 24.7 -12.98 25.05 -12.86 ;
      RECT 24.7 -9.75 25.05 -9.63 ;
      RECT 24.7 -6.52 25.05 -6.4 ;
      RECT 24.7 -3.29 25.05 -3.17 ;
      RECT 24.7 -0.06 25.05 0.06 ;
      RECT 24.815 -56.495 24.915 -55.535 ;
      RECT 24.815 2.175 24.915 3.135 ;
      RECT 24.715 -61.875 24.815 -61.405 ;
      RECT 24.215 -48.51 24.565 -48.39 ;
      RECT 24.215 -45.28 24.565 -45.16 ;
      RECT 24.215 -42.05 24.565 -41.93 ;
      RECT 24.215 -38.82 24.565 -38.7 ;
      RECT 24.215 -35.59 24.565 -35.47 ;
      RECT 24.215 -32.36 24.565 -32.24 ;
      RECT 24.215 -29.13 24.565 -29.01 ;
      RECT 24.215 -25.9 24.565 -25.78 ;
      RECT 24.215 -22.67 24.565 -22.55 ;
      RECT 24.215 -19.44 24.565 -19.32 ;
      RECT 24.215 -16.21 24.565 -16.09 ;
      RECT 24.215 -12.98 24.565 -12.86 ;
      RECT 24.215 -9.75 24.565 -9.63 ;
      RECT 24.215 -6.52 24.565 -6.4 ;
      RECT 24.215 -3.29 24.565 -3.17 ;
      RECT 24.215 -0.06 24.565 0.06 ;
      RECT 24.35 -59.055 24.5 -58.765 ;
      RECT 24.385 -56.495 24.485 -55.535 ;
      RECT 24.385 2.175 24.485 3.135 ;
      RECT 24.365 -60.51 24.465 -59.97 ;
      RECT 24.125 -61.875 24.225 -61.405 ;
      RECT 24.125 -56.495 24.225 -55.535 ;
      RECT 23.875 -53.265 23.975 -52.305 ;
      RECT 23.5 -48.51 23.85 -48.39 ;
      RECT 23.5 -45.28 23.85 -45.16 ;
      RECT 23.5 -42.05 23.85 -41.93 ;
      RECT 23.5 -38.82 23.85 -38.7 ;
      RECT 23.5 -35.59 23.85 -35.47 ;
      RECT 23.5 -32.36 23.85 -32.24 ;
      RECT 23.5 -29.13 23.85 -29.01 ;
      RECT 23.5 -25.9 23.85 -25.78 ;
      RECT 23.5 -22.67 23.85 -22.55 ;
      RECT 23.5 -19.44 23.85 -19.32 ;
      RECT 23.5 -16.21 23.85 -16.09 ;
      RECT 23.5 -12.98 23.85 -12.86 ;
      RECT 23.5 -9.75 23.85 -9.63 ;
      RECT 23.5 -6.52 23.85 -6.4 ;
      RECT 23.5 -3.29 23.85 -3.17 ;
      RECT 23.5 -0.06 23.85 0.06 ;
      RECT 23.615 -53.265 23.715 -52.305 ;
      RECT 23.615 2.175 23.715 3.135 ;
      RECT 23.325 -60.575 23.425 -60.095 ;
      RECT 23.325 -59.085 23.425 -58.615 ;
      RECT 23.015 -48.51 23.365 -48.39 ;
      RECT 23.015 -45.28 23.365 -45.16 ;
      RECT 23.015 -42.05 23.365 -41.93 ;
      RECT 23.015 -38.82 23.365 -38.7 ;
      RECT 23.015 -35.59 23.365 -35.47 ;
      RECT 23.015 -32.36 23.365 -32.24 ;
      RECT 23.015 -29.13 23.365 -29.01 ;
      RECT 23.015 -25.9 23.365 -25.78 ;
      RECT 23.015 -22.67 23.365 -22.55 ;
      RECT 23.015 -19.44 23.365 -19.32 ;
      RECT 23.015 -16.21 23.365 -16.09 ;
      RECT 23.015 -12.98 23.365 -12.86 ;
      RECT 23.015 -9.75 23.365 -9.63 ;
      RECT 23.015 -6.52 23.365 -6.4 ;
      RECT 23.015 -3.29 23.365 -3.17 ;
      RECT 23.015 -0.06 23.365 0.06 ;
      RECT 23.185 -53.265 23.285 -52.305 ;
      RECT 23.185 2.175 23.285 3.135 ;
      RECT 19.285 -56.975 23.065 -56.855 ;
      RECT 22.925 -53.265 23.025 -52.305 ;
      RECT 22.735 -59.07 22.855 -58.69 ;
      RECT 22.735 -60.565 22.835 -60.095 ;
      RECT 22.675 -53.265 22.775 -52.305 ;
      RECT 22.3 -48.51 22.65 -48.39 ;
      RECT 22.3 -45.28 22.65 -45.16 ;
      RECT 22.3 -42.05 22.65 -41.93 ;
      RECT 22.3 -38.82 22.65 -38.7 ;
      RECT 22.3 -35.59 22.65 -35.47 ;
      RECT 22.3 -32.36 22.65 -32.24 ;
      RECT 22.3 -29.13 22.65 -29.01 ;
      RECT 22.3 -25.9 22.65 -25.78 ;
      RECT 22.3 -22.67 22.65 -22.55 ;
      RECT 22.3 -19.44 22.65 -19.32 ;
      RECT 22.3 -16.21 22.65 -16.09 ;
      RECT 22.3 -12.98 22.65 -12.86 ;
      RECT 22.3 -9.75 22.65 -9.63 ;
      RECT 22.3 -6.52 22.65 -6.4 ;
      RECT 22.3 -3.29 22.65 -3.17 ;
      RECT 22.3 -0.06 22.65 0.06 ;
      RECT 22.415 -53.265 22.515 -52.305 ;
      RECT 22.415 2.175 22.515 3.135 ;
      RECT 22.145 -57.915 22.28 -57.595 ;
      RECT 21.815 -48.51 22.165 -48.39 ;
      RECT 21.815 -45.28 22.165 -45.16 ;
      RECT 21.815 -42.05 22.165 -41.93 ;
      RECT 21.815 -38.82 22.165 -38.7 ;
      RECT 21.815 -35.59 22.165 -35.47 ;
      RECT 21.815 -32.36 22.165 -32.24 ;
      RECT 21.815 -29.13 22.165 -29.01 ;
      RECT 21.815 -25.9 22.165 -25.78 ;
      RECT 21.815 -22.67 22.165 -22.55 ;
      RECT 21.815 -19.44 22.165 -19.32 ;
      RECT 21.815 -16.21 22.165 -16.09 ;
      RECT 21.815 -12.98 22.165 -12.86 ;
      RECT 21.815 -9.75 22.165 -9.63 ;
      RECT 21.815 -6.52 22.165 -6.4 ;
      RECT 21.815 -3.29 22.165 -3.17 ;
      RECT 21.815 -0.06 22.165 0.06 ;
      RECT 21.985 -53.265 22.085 -52.305 ;
      RECT 21.985 2.175 22.085 3.135 ;
      RECT 21.81 -57.915 21.955 -57.595 ;
      RECT 21.725 -53.265 21.825 -52.305 ;
      RECT 21.475 -56.495 21.575 -55.535 ;
      RECT 21.1 -48.51 21.45 -48.39 ;
      RECT 21.1 -45.28 21.45 -45.16 ;
      RECT 21.1 -42.05 21.45 -41.93 ;
      RECT 21.1 -38.82 21.45 -38.7 ;
      RECT 21.1 -35.59 21.45 -35.47 ;
      RECT 21.1 -32.36 21.45 -32.24 ;
      RECT 21.1 -29.13 21.45 -29.01 ;
      RECT 21.1 -25.9 21.45 -25.78 ;
      RECT 21.1 -22.67 21.45 -22.55 ;
      RECT 21.1 -19.44 21.45 -19.32 ;
      RECT 21.1 -16.21 21.45 -16.09 ;
      RECT 21.1 -12.98 21.45 -12.86 ;
      RECT 21.1 -9.75 21.45 -9.63 ;
      RECT 21.1 -6.52 21.45 -6.4 ;
      RECT 21.1 -3.29 21.45 -3.17 ;
      RECT 21.1 -0.06 21.45 0.06 ;
      RECT 21.305 -60.575 21.405 -60.095 ;
      RECT 21.305 -59.085 21.405 -58.615 ;
      RECT 21.215 -56.495 21.315 -55.535 ;
      RECT 21.215 2.175 21.315 3.135 ;
      RECT 20.615 -48.51 20.965 -48.39 ;
      RECT 20.615 -45.28 20.965 -45.16 ;
      RECT 20.615 -42.05 20.965 -41.93 ;
      RECT 20.615 -38.82 20.965 -38.7 ;
      RECT 20.615 -35.59 20.965 -35.47 ;
      RECT 20.615 -32.36 20.965 -32.24 ;
      RECT 20.615 -29.13 20.965 -29.01 ;
      RECT 20.615 -25.9 20.965 -25.78 ;
      RECT 20.615 -22.67 20.965 -22.55 ;
      RECT 20.615 -19.44 20.965 -19.32 ;
      RECT 20.615 -16.21 20.965 -16.09 ;
      RECT 20.615 -12.98 20.965 -12.86 ;
      RECT 20.615 -9.75 20.965 -9.63 ;
      RECT 20.615 -6.52 20.965 -6.4 ;
      RECT 20.615 -3.29 20.965 -3.17 ;
      RECT 20.615 -0.06 20.965 0.06 ;
      RECT 20.785 -56.495 20.885 -55.535 ;
      RECT 20.785 2.175 20.885 3.135 ;
      RECT 20.68 -59.085 20.85 -58.705 ;
      RECT 20.715 -60.565 20.815 -60.095 ;
      RECT 20.525 -56.495 20.625 -55.535 ;
      RECT 20.275 -56.495 20.375 -55.535 ;
      RECT 19.9 -48.51 20.25 -48.39 ;
      RECT 19.9 -45.28 20.25 -45.16 ;
      RECT 19.9 -42.05 20.25 -41.93 ;
      RECT 19.9 -38.82 20.25 -38.7 ;
      RECT 19.9 -35.59 20.25 -35.47 ;
      RECT 19.9 -32.36 20.25 -32.24 ;
      RECT 19.9 -29.13 20.25 -29.01 ;
      RECT 19.9 -25.9 20.25 -25.78 ;
      RECT 19.9 -22.67 20.25 -22.55 ;
      RECT 19.9 -19.44 20.25 -19.32 ;
      RECT 19.9 -16.21 20.25 -16.09 ;
      RECT 19.9 -12.98 20.25 -12.86 ;
      RECT 19.9 -9.75 20.25 -9.63 ;
      RECT 19.9 -6.52 20.25 -6.4 ;
      RECT 19.9 -3.29 20.25 -3.17 ;
      RECT 19.9 -0.06 20.25 0.06 ;
      RECT 20.015 -56.495 20.115 -55.535 ;
      RECT 20.015 2.175 20.115 3.135 ;
      RECT 19.915 -61.875 20.015 -61.405 ;
      RECT 19.415 -48.51 19.765 -48.39 ;
      RECT 19.415 -45.28 19.765 -45.16 ;
      RECT 19.415 -42.05 19.765 -41.93 ;
      RECT 19.415 -38.82 19.765 -38.7 ;
      RECT 19.415 -35.59 19.765 -35.47 ;
      RECT 19.415 -32.36 19.765 -32.24 ;
      RECT 19.415 -29.13 19.765 -29.01 ;
      RECT 19.415 -25.9 19.765 -25.78 ;
      RECT 19.415 -22.67 19.765 -22.55 ;
      RECT 19.415 -19.44 19.765 -19.32 ;
      RECT 19.415 -16.21 19.765 -16.09 ;
      RECT 19.415 -12.98 19.765 -12.86 ;
      RECT 19.415 -9.75 19.765 -9.63 ;
      RECT 19.415 -6.52 19.765 -6.4 ;
      RECT 19.415 -3.29 19.765 -3.17 ;
      RECT 19.415 -0.06 19.765 0.06 ;
      RECT 19.55 -59.055 19.7 -58.765 ;
      RECT 19.585 -56.495 19.685 -55.535 ;
      RECT 19.585 2.175 19.685 3.135 ;
      RECT 19.565 -60.51 19.665 -59.97 ;
      RECT 19.325 -61.875 19.425 -61.405 ;
      RECT 19.325 -56.495 19.425 -55.535 ;
      RECT 19.075 -53.265 19.175 -52.305 ;
      RECT 18.7 -48.51 19.05 -48.39 ;
      RECT 18.7 -45.28 19.05 -45.16 ;
      RECT 18.7 -42.05 19.05 -41.93 ;
      RECT 18.7 -38.82 19.05 -38.7 ;
      RECT 18.7 -35.59 19.05 -35.47 ;
      RECT 18.7 -32.36 19.05 -32.24 ;
      RECT 18.7 -29.13 19.05 -29.01 ;
      RECT 18.7 -25.9 19.05 -25.78 ;
      RECT 18.7 -22.67 19.05 -22.55 ;
      RECT 18.7 -19.44 19.05 -19.32 ;
      RECT 18.7 -16.21 19.05 -16.09 ;
      RECT 18.7 -12.98 19.05 -12.86 ;
      RECT 18.7 -9.75 19.05 -9.63 ;
      RECT 18.7 -6.52 19.05 -6.4 ;
      RECT 18.7 -3.29 19.05 -3.17 ;
      RECT 18.7 -0.06 19.05 0.06 ;
      RECT 18.815 -53.265 18.915 -52.305 ;
      RECT 18.815 2.175 18.915 3.135 ;
      RECT 18.525 -60.575 18.625 -60.095 ;
      RECT 18.525 -59.085 18.625 -58.615 ;
      RECT 18.215 -48.51 18.565 -48.39 ;
      RECT 18.215 -45.28 18.565 -45.16 ;
      RECT 18.215 -42.05 18.565 -41.93 ;
      RECT 18.215 -38.82 18.565 -38.7 ;
      RECT 18.215 -35.59 18.565 -35.47 ;
      RECT 18.215 -32.36 18.565 -32.24 ;
      RECT 18.215 -29.13 18.565 -29.01 ;
      RECT 18.215 -25.9 18.565 -25.78 ;
      RECT 18.215 -22.67 18.565 -22.55 ;
      RECT 18.215 -19.44 18.565 -19.32 ;
      RECT 18.215 -16.21 18.565 -16.09 ;
      RECT 18.215 -12.98 18.565 -12.86 ;
      RECT 18.215 -9.75 18.565 -9.63 ;
      RECT 18.215 -6.52 18.565 -6.4 ;
      RECT 18.215 -3.29 18.565 -3.17 ;
      RECT 18.215 -0.06 18.565 0.06 ;
      RECT 18.385 -53.265 18.485 -52.305 ;
      RECT 18.385 2.175 18.485 3.135 ;
      RECT 14.485 -56.975 18.265 -56.855 ;
      RECT 18.125 -53.265 18.225 -52.305 ;
      RECT 17.935 -59.07 18.055 -58.69 ;
      RECT 17.935 -60.565 18.035 -60.095 ;
      RECT 17.875 -53.265 17.975 -52.305 ;
      RECT 17.5 -48.51 17.85 -48.39 ;
      RECT 17.5 -45.28 17.85 -45.16 ;
      RECT 17.5 -42.05 17.85 -41.93 ;
      RECT 17.5 -38.82 17.85 -38.7 ;
      RECT 17.5 -35.59 17.85 -35.47 ;
      RECT 17.5 -32.36 17.85 -32.24 ;
      RECT 17.5 -29.13 17.85 -29.01 ;
      RECT 17.5 -25.9 17.85 -25.78 ;
      RECT 17.5 -22.67 17.85 -22.55 ;
      RECT 17.5 -19.44 17.85 -19.32 ;
      RECT 17.5 -16.21 17.85 -16.09 ;
      RECT 17.5 -12.98 17.85 -12.86 ;
      RECT 17.5 -9.75 17.85 -9.63 ;
      RECT 17.5 -6.52 17.85 -6.4 ;
      RECT 17.5 -3.29 17.85 -3.17 ;
      RECT 17.5 -0.06 17.85 0.06 ;
      RECT 17.615 -53.265 17.715 -52.305 ;
      RECT 17.615 2.175 17.715 3.135 ;
      RECT 17.345 -57.915 17.48 -57.595 ;
      RECT 17.015 -48.51 17.365 -48.39 ;
      RECT 17.015 -45.28 17.365 -45.16 ;
      RECT 17.015 -42.05 17.365 -41.93 ;
      RECT 17.015 -38.82 17.365 -38.7 ;
      RECT 17.015 -35.59 17.365 -35.47 ;
      RECT 17.015 -32.36 17.365 -32.24 ;
      RECT 17.015 -29.13 17.365 -29.01 ;
      RECT 17.015 -25.9 17.365 -25.78 ;
      RECT 17.015 -22.67 17.365 -22.55 ;
      RECT 17.015 -19.44 17.365 -19.32 ;
      RECT 17.015 -16.21 17.365 -16.09 ;
      RECT 17.015 -12.98 17.365 -12.86 ;
      RECT 17.015 -9.75 17.365 -9.63 ;
      RECT 17.015 -6.52 17.365 -6.4 ;
      RECT 17.015 -3.29 17.365 -3.17 ;
      RECT 17.015 -0.06 17.365 0.06 ;
      RECT 17.185 -53.265 17.285 -52.305 ;
      RECT 17.185 2.175 17.285 3.135 ;
      RECT 17.01 -57.915 17.155 -57.595 ;
      RECT 16.925 -53.265 17.025 -52.305 ;
      RECT 16.675 -56.495 16.775 -55.535 ;
      RECT 16.3 -48.51 16.65 -48.39 ;
      RECT 16.3 -45.28 16.65 -45.16 ;
      RECT 16.3 -42.05 16.65 -41.93 ;
      RECT 16.3 -38.82 16.65 -38.7 ;
      RECT 16.3 -35.59 16.65 -35.47 ;
      RECT 16.3 -32.36 16.65 -32.24 ;
      RECT 16.3 -29.13 16.65 -29.01 ;
      RECT 16.3 -25.9 16.65 -25.78 ;
      RECT 16.3 -22.67 16.65 -22.55 ;
      RECT 16.3 -19.44 16.65 -19.32 ;
      RECT 16.3 -16.21 16.65 -16.09 ;
      RECT 16.3 -12.98 16.65 -12.86 ;
      RECT 16.3 -9.75 16.65 -9.63 ;
      RECT 16.3 -6.52 16.65 -6.4 ;
      RECT 16.3 -3.29 16.65 -3.17 ;
      RECT 16.3 -0.06 16.65 0.06 ;
      RECT 16.505 -60.575 16.605 -60.095 ;
      RECT 16.505 -59.085 16.605 -58.615 ;
      RECT 16.415 -56.495 16.515 -55.535 ;
      RECT 16.415 2.175 16.515 3.135 ;
      RECT 15.815 -48.51 16.165 -48.39 ;
      RECT 15.815 -45.28 16.165 -45.16 ;
      RECT 15.815 -42.05 16.165 -41.93 ;
      RECT 15.815 -38.82 16.165 -38.7 ;
      RECT 15.815 -35.59 16.165 -35.47 ;
      RECT 15.815 -32.36 16.165 -32.24 ;
      RECT 15.815 -29.13 16.165 -29.01 ;
      RECT 15.815 -25.9 16.165 -25.78 ;
      RECT 15.815 -22.67 16.165 -22.55 ;
      RECT 15.815 -19.44 16.165 -19.32 ;
      RECT 15.815 -16.21 16.165 -16.09 ;
      RECT 15.815 -12.98 16.165 -12.86 ;
      RECT 15.815 -9.75 16.165 -9.63 ;
      RECT 15.815 -6.52 16.165 -6.4 ;
      RECT 15.815 -3.29 16.165 -3.17 ;
      RECT 15.815 -0.06 16.165 0.06 ;
      RECT 15.985 -56.495 16.085 -55.535 ;
      RECT 15.985 2.175 16.085 3.135 ;
      RECT 15.88 -59.085 16.05 -58.705 ;
      RECT 15.915 -60.565 16.015 -60.095 ;
      RECT 15.725 -56.495 15.825 -55.535 ;
      RECT 15.475 -56.495 15.575 -55.535 ;
      RECT 15.1 -48.51 15.45 -48.39 ;
      RECT 15.1 -45.28 15.45 -45.16 ;
      RECT 15.1 -42.05 15.45 -41.93 ;
      RECT 15.1 -38.82 15.45 -38.7 ;
      RECT 15.1 -35.59 15.45 -35.47 ;
      RECT 15.1 -32.36 15.45 -32.24 ;
      RECT 15.1 -29.13 15.45 -29.01 ;
      RECT 15.1 -25.9 15.45 -25.78 ;
      RECT 15.1 -22.67 15.45 -22.55 ;
      RECT 15.1 -19.44 15.45 -19.32 ;
      RECT 15.1 -16.21 15.45 -16.09 ;
      RECT 15.1 -12.98 15.45 -12.86 ;
      RECT 15.1 -9.75 15.45 -9.63 ;
      RECT 15.1 -6.52 15.45 -6.4 ;
      RECT 15.1 -3.29 15.45 -3.17 ;
      RECT 15.1 -0.06 15.45 0.06 ;
      RECT 15.215 -56.495 15.315 -55.535 ;
      RECT 15.215 2.175 15.315 3.135 ;
      RECT 15.115 -61.875 15.215 -61.405 ;
      RECT 14.615 -48.51 14.965 -48.39 ;
      RECT 14.615 -45.28 14.965 -45.16 ;
      RECT 14.615 -42.05 14.965 -41.93 ;
      RECT 14.615 -38.82 14.965 -38.7 ;
      RECT 14.615 -35.59 14.965 -35.47 ;
      RECT 14.615 -32.36 14.965 -32.24 ;
      RECT 14.615 -29.13 14.965 -29.01 ;
      RECT 14.615 -25.9 14.965 -25.78 ;
      RECT 14.615 -22.67 14.965 -22.55 ;
      RECT 14.615 -19.44 14.965 -19.32 ;
      RECT 14.615 -16.21 14.965 -16.09 ;
      RECT 14.615 -12.98 14.965 -12.86 ;
      RECT 14.615 -9.75 14.965 -9.63 ;
      RECT 14.615 -6.52 14.965 -6.4 ;
      RECT 14.615 -3.29 14.965 -3.17 ;
      RECT 14.615 -0.06 14.965 0.06 ;
      RECT 14.75 -59.055 14.9 -58.765 ;
      RECT 14.785 -56.495 14.885 -55.535 ;
      RECT 14.785 2.175 14.885 3.135 ;
      RECT 14.765 -60.51 14.865 -59.97 ;
      RECT 14.525 -61.875 14.625 -61.405 ;
      RECT 14.525 -56.495 14.625 -55.535 ;
      RECT 14.275 -53.265 14.375 -52.305 ;
      RECT 13.9 -48.51 14.25 -48.39 ;
      RECT 13.9 -45.28 14.25 -45.16 ;
      RECT 13.9 -42.05 14.25 -41.93 ;
      RECT 13.9 -38.82 14.25 -38.7 ;
      RECT 13.9 -35.59 14.25 -35.47 ;
      RECT 13.9 -32.36 14.25 -32.24 ;
      RECT 13.9 -29.13 14.25 -29.01 ;
      RECT 13.9 -25.9 14.25 -25.78 ;
      RECT 13.9 -22.67 14.25 -22.55 ;
      RECT 13.9 -19.44 14.25 -19.32 ;
      RECT 13.9 -16.21 14.25 -16.09 ;
      RECT 13.9 -12.98 14.25 -12.86 ;
      RECT 13.9 -9.75 14.25 -9.63 ;
      RECT 13.9 -6.52 14.25 -6.4 ;
      RECT 13.9 -3.29 14.25 -3.17 ;
      RECT 13.9 -0.06 14.25 0.06 ;
      RECT 14.015 -53.265 14.115 -52.305 ;
      RECT 14.015 2.175 14.115 3.135 ;
      RECT 13.725 -60.575 13.825 -60.095 ;
      RECT 13.725 -59.085 13.825 -58.615 ;
      RECT 13.415 -48.51 13.765 -48.39 ;
      RECT 13.415 -45.28 13.765 -45.16 ;
      RECT 13.415 -42.05 13.765 -41.93 ;
      RECT 13.415 -38.82 13.765 -38.7 ;
      RECT 13.415 -35.59 13.765 -35.47 ;
      RECT 13.415 -32.36 13.765 -32.24 ;
      RECT 13.415 -29.13 13.765 -29.01 ;
      RECT 13.415 -25.9 13.765 -25.78 ;
      RECT 13.415 -22.67 13.765 -22.55 ;
      RECT 13.415 -19.44 13.765 -19.32 ;
      RECT 13.415 -16.21 13.765 -16.09 ;
      RECT 13.415 -12.98 13.765 -12.86 ;
      RECT 13.415 -9.75 13.765 -9.63 ;
      RECT 13.415 -6.52 13.765 -6.4 ;
      RECT 13.415 -3.29 13.765 -3.17 ;
      RECT 13.415 -0.06 13.765 0.06 ;
      RECT 13.585 -53.265 13.685 -52.305 ;
      RECT 13.585 2.175 13.685 3.135 ;
      RECT 9.685 -56.975 13.465 -56.855 ;
      RECT 13.325 -53.265 13.425 -52.305 ;
      RECT 13.135 -59.07 13.255 -58.69 ;
      RECT 13.135 -60.565 13.235 -60.095 ;
      RECT 13.075 -53.265 13.175 -52.305 ;
      RECT 12.7 -48.51 13.05 -48.39 ;
      RECT 12.7 -45.28 13.05 -45.16 ;
      RECT 12.7 -42.05 13.05 -41.93 ;
      RECT 12.7 -38.82 13.05 -38.7 ;
      RECT 12.7 -35.59 13.05 -35.47 ;
      RECT 12.7 -32.36 13.05 -32.24 ;
      RECT 12.7 -29.13 13.05 -29.01 ;
      RECT 12.7 -25.9 13.05 -25.78 ;
      RECT 12.7 -22.67 13.05 -22.55 ;
      RECT 12.7 -19.44 13.05 -19.32 ;
      RECT 12.7 -16.21 13.05 -16.09 ;
      RECT 12.7 -12.98 13.05 -12.86 ;
      RECT 12.7 -9.75 13.05 -9.63 ;
      RECT 12.7 -6.52 13.05 -6.4 ;
      RECT 12.7 -3.29 13.05 -3.17 ;
      RECT 12.7 -0.06 13.05 0.06 ;
      RECT 12.815 -53.265 12.915 -52.305 ;
      RECT 12.815 2.175 12.915 3.135 ;
      RECT 12.545 -57.915 12.68 -57.595 ;
      RECT 12.215 -48.51 12.565 -48.39 ;
      RECT 12.215 -45.28 12.565 -45.16 ;
      RECT 12.215 -42.05 12.565 -41.93 ;
      RECT 12.215 -38.82 12.565 -38.7 ;
      RECT 12.215 -35.59 12.565 -35.47 ;
      RECT 12.215 -32.36 12.565 -32.24 ;
      RECT 12.215 -29.13 12.565 -29.01 ;
      RECT 12.215 -25.9 12.565 -25.78 ;
      RECT 12.215 -22.67 12.565 -22.55 ;
      RECT 12.215 -19.44 12.565 -19.32 ;
      RECT 12.215 -16.21 12.565 -16.09 ;
      RECT 12.215 -12.98 12.565 -12.86 ;
      RECT 12.215 -9.75 12.565 -9.63 ;
      RECT 12.215 -6.52 12.565 -6.4 ;
      RECT 12.215 -3.29 12.565 -3.17 ;
      RECT 12.215 -0.06 12.565 0.06 ;
      RECT 12.385 -53.265 12.485 -52.305 ;
      RECT 12.385 2.175 12.485 3.135 ;
      RECT 12.21 -57.915 12.355 -57.595 ;
      RECT 12.125 -53.265 12.225 -52.305 ;
      RECT 11.875 -56.495 11.975 -55.535 ;
      RECT 11.5 -48.51 11.85 -48.39 ;
      RECT 11.5 -45.28 11.85 -45.16 ;
      RECT 11.5 -42.05 11.85 -41.93 ;
      RECT 11.5 -38.82 11.85 -38.7 ;
      RECT 11.5 -35.59 11.85 -35.47 ;
      RECT 11.5 -32.36 11.85 -32.24 ;
      RECT 11.5 -29.13 11.85 -29.01 ;
      RECT 11.5 -25.9 11.85 -25.78 ;
      RECT 11.5 -22.67 11.85 -22.55 ;
      RECT 11.5 -19.44 11.85 -19.32 ;
      RECT 11.5 -16.21 11.85 -16.09 ;
      RECT 11.5 -12.98 11.85 -12.86 ;
      RECT 11.5 -9.75 11.85 -9.63 ;
      RECT 11.5 -6.52 11.85 -6.4 ;
      RECT 11.5 -3.29 11.85 -3.17 ;
      RECT 11.5 -0.06 11.85 0.06 ;
      RECT 11.705 -60.575 11.805 -60.095 ;
      RECT 11.705 -59.085 11.805 -58.615 ;
      RECT 11.615 -56.495 11.715 -55.535 ;
      RECT 11.615 2.175 11.715 3.135 ;
      RECT 11.015 -48.51 11.365 -48.39 ;
      RECT 11.015 -45.28 11.365 -45.16 ;
      RECT 11.015 -42.05 11.365 -41.93 ;
      RECT 11.015 -38.82 11.365 -38.7 ;
      RECT 11.015 -35.59 11.365 -35.47 ;
      RECT 11.015 -32.36 11.365 -32.24 ;
      RECT 11.015 -29.13 11.365 -29.01 ;
      RECT 11.015 -25.9 11.365 -25.78 ;
      RECT 11.015 -22.67 11.365 -22.55 ;
      RECT 11.015 -19.44 11.365 -19.32 ;
      RECT 11.015 -16.21 11.365 -16.09 ;
      RECT 11.015 -12.98 11.365 -12.86 ;
      RECT 11.015 -9.75 11.365 -9.63 ;
      RECT 11.015 -6.52 11.365 -6.4 ;
      RECT 11.015 -3.29 11.365 -3.17 ;
      RECT 11.015 -0.06 11.365 0.06 ;
      RECT 11.185 -56.495 11.285 -55.535 ;
      RECT 11.185 2.175 11.285 3.135 ;
      RECT 11.08 -59.085 11.25 -58.705 ;
      RECT 11.115 -60.565 11.215 -60.095 ;
      RECT 10.925 -56.495 11.025 -55.535 ;
      RECT 10.675 -56.495 10.775 -55.535 ;
      RECT 10.3 -48.51 10.65 -48.39 ;
      RECT 10.3 -45.28 10.65 -45.16 ;
      RECT 10.3 -42.05 10.65 -41.93 ;
      RECT 10.3 -38.82 10.65 -38.7 ;
      RECT 10.3 -35.59 10.65 -35.47 ;
      RECT 10.3 -32.36 10.65 -32.24 ;
      RECT 10.3 -29.13 10.65 -29.01 ;
      RECT 10.3 -25.9 10.65 -25.78 ;
      RECT 10.3 -22.67 10.65 -22.55 ;
      RECT 10.3 -19.44 10.65 -19.32 ;
      RECT 10.3 -16.21 10.65 -16.09 ;
      RECT 10.3 -12.98 10.65 -12.86 ;
      RECT 10.3 -9.75 10.65 -9.63 ;
      RECT 10.3 -6.52 10.65 -6.4 ;
      RECT 10.3 -3.29 10.65 -3.17 ;
      RECT 10.3 -0.06 10.65 0.06 ;
      RECT 10.415 -56.495 10.515 -55.535 ;
      RECT 10.415 2.175 10.515 3.135 ;
      RECT 10.315 -61.875 10.415 -61.405 ;
      RECT 9.815 -48.51 10.165 -48.39 ;
      RECT 9.815 -45.28 10.165 -45.16 ;
      RECT 9.815 -42.05 10.165 -41.93 ;
      RECT 9.815 -38.82 10.165 -38.7 ;
      RECT 9.815 -35.59 10.165 -35.47 ;
      RECT 9.815 -32.36 10.165 -32.24 ;
      RECT 9.815 -29.13 10.165 -29.01 ;
      RECT 9.815 -25.9 10.165 -25.78 ;
      RECT 9.815 -22.67 10.165 -22.55 ;
      RECT 9.815 -19.44 10.165 -19.32 ;
      RECT 9.815 -16.21 10.165 -16.09 ;
      RECT 9.815 -12.98 10.165 -12.86 ;
      RECT 9.815 -9.75 10.165 -9.63 ;
      RECT 9.815 -6.52 10.165 -6.4 ;
      RECT 9.815 -3.29 10.165 -3.17 ;
      RECT 9.815 -0.06 10.165 0.06 ;
      RECT 9.95 -59.055 10.1 -58.765 ;
      RECT 9.985 -56.495 10.085 -55.535 ;
      RECT 9.985 2.175 10.085 3.135 ;
      RECT 9.965 -60.51 10.065 -59.97 ;
      RECT 9.725 -61.875 9.825 -61.405 ;
      RECT 9.725 -56.495 9.825 -55.535 ;
      RECT 9.475 -53.265 9.575 -52.305 ;
      RECT 9.1 -48.51 9.45 -48.39 ;
      RECT 9.1 -45.28 9.45 -45.16 ;
      RECT 9.1 -42.05 9.45 -41.93 ;
      RECT 9.1 -38.82 9.45 -38.7 ;
      RECT 9.1 -35.59 9.45 -35.47 ;
      RECT 9.1 -32.36 9.45 -32.24 ;
      RECT 9.1 -29.13 9.45 -29.01 ;
      RECT 9.1 -25.9 9.45 -25.78 ;
      RECT 9.1 -22.67 9.45 -22.55 ;
      RECT 9.1 -19.44 9.45 -19.32 ;
      RECT 9.1 -16.21 9.45 -16.09 ;
      RECT 9.1 -12.98 9.45 -12.86 ;
      RECT 9.1 -9.75 9.45 -9.63 ;
      RECT 9.1 -6.52 9.45 -6.4 ;
      RECT 9.1 -3.29 9.45 -3.17 ;
      RECT 9.1 -0.06 9.45 0.06 ;
      RECT 9.215 -53.265 9.315 -52.305 ;
      RECT 9.215 2.175 9.315 3.135 ;
      RECT 8.925 -60.575 9.025 -60.095 ;
      RECT 8.925 -59.085 9.025 -58.615 ;
      RECT 8.615 -48.51 8.965 -48.39 ;
      RECT 8.615 -45.28 8.965 -45.16 ;
      RECT 8.615 -42.05 8.965 -41.93 ;
      RECT 8.615 -38.82 8.965 -38.7 ;
      RECT 8.615 -35.59 8.965 -35.47 ;
      RECT 8.615 -32.36 8.965 -32.24 ;
      RECT 8.615 -29.13 8.965 -29.01 ;
      RECT 8.615 -25.9 8.965 -25.78 ;
      RECT 8.615 -22.67 8.965 -22.55 ;
      RECT 8.615 -19.44 8.965 -19.32 ;
      RECT 8.615 -16.21 8.965 -16.09 ;
      RECT 8.615 -12.98 8.965 -12.86 ;
      RECT 8.615 -9.75 8.965 -9.63 ;
      RECT 8.615 -6.52 8.965 -6.4 ;
      RECT 8.615 -3.29 8.965 -3.17 ;
      RECT 8.615 -0.06 8.965 0.06 ;
      RECT 8.785 -53.265 8.885 -52.305 ;
      RECT 8.785 2.175 8.885 3.135 ;
      RECT 4.885 -56.975 8.665 -56.855 ;
      RECT 8.525 -53.265 8.625 -52.305 ;
      RECT 8.335 -59.07 8.455 -58.69 ;
      RECT 8.335 -60.565 8.435 -60.095 ;
      RECT 8.275 -53.265 8.375 -52.305 ;
      RECT 7.9 -48.51 8.25 -48.39 ;
      RECT 7.9 -45.28 8.25 -45.16 ;
      RECT 7.9 -42.05 8.25 -41.93 ;
      RECT 7.9 -38.82 8.25 -38.7 ;
      RECT 7.9 -35.59 8.25 -35.47 ;
      RECT 7.9 -32.36 8.25 -32.24 ;
      RECT 7.9 -29.13 8.25 -29.01 ;
      RECT 7.9 -25.9 8.25 -25.78 ;
      RECT 7.9 -22.67 8.25 -22.55 ;
      RECT 7.9 -19.44 8.25 -19.32 ;
      RECT 7.9 -16.21 8.25 -16.09 ;
      RECT 7.9 -12.98 8.25 -12.86 ;
      RECT 7.9 -9.75 8.25 -9.63 ;
      RECT 7.9 -6.52 8.25 -6.4 ;
      RECT 7.9 -3.29 8.25 -3.17 ;
      RECT 7.9 -0.06 8.25 0.06 ;
      RECT 8.015 -53.265 8.115 -52.305 ;
      RECT 8.015 2.175 8.115 3.135 ;
      RECT 7.745 -57.915 7.88 -57.595 ;
      RECT 7.415 -48.51 7.765 -48.39 ;
      RECT 7.415 -45.28 7.765 -45.16 ;
      RECT 7.415 -42.05 7.765 -41.93 ;
      RECT 7.415 -38.82 7.765 -38.7 ;
      RECT 7.415 -35.59 7.765 -35.47 ;
      RECT 7.415 -32.36 7.765 -32.24 ;
      RECT 7.415 -29.13 7.765 -29.01 ;
      RECT 7.415 -25.9 7.765 -25.78 ;
      RECT 7.415 -22.67 7.765 -22.55 ;
      RECT 7.415 -19.44 7.765 -19.32 ;
      RECT 7.415 -16.21 7.765 -16.09 ;
      RECT 7.415 -12.98 7.765 -12.86 ;
      RECT 7.415 -9.75 7.765 -9.63 ;
      RECT 7.415 -6.52 7.765 -6.4 ;
      RECT 7.415 -3.29 7.765 -3.17 ;
      RECT 7.415 -0.06 7.765 0.06 ;
      RECT 7.585 -53.265 7.685 -52.305 ;
      RECT 7.585 2.175 7.685 3.135 ;
      RECT 7.41 -57.915 7.555 -57.595 ;
      RECT 7.325 -53.265 7.425 -52.305 ;
      RECT 7.075 -56.495 7.175 -55.535 ;
      RECT 6.7 -48.51 7.05 -48.39 ;
      RECT 6.7 -45.28 7.05 -45.16 ;
      RECT 6.7 -42.05 7.05 -41.93 ;
      RECT 6.7 -38.82 7.05 -38.7 ;
      RECT 6.7 -35.59 7.05 -35.47 ;
      RECT 6.7 -32.36 7.05 -32.24 ;
      RECT 6.7 -29.13 7.05 -29.01 ;
      RECT 6.7 -25.9 7.05 -25.78 ;
      RECT 6.7 -22.67 7.05 -22.55 ;
      RECT 6.7 -19.44 7.05 -19.32 ;
      RECT 6.7 -16.21 7.05 -16.09 ;
      RECT 6.7 -12.98 7.05 -12.86 ;
      RECT 6.7 -9.75 7.05 -9.63 ;
      RECT 6.7 -6.52 7.05 -6.4 ;
      RECT 6.7 -3.29 7.05 -3.17 ;
      RECT 6.7 -0.06 7.05 0.06 ;
      RECT 6.905 -60.575 7.005 -60.095 ;
      RECT 6.905 -59.085 7.005 -58.615 ;
      RECT 6.815 -56.495 6.915 -55.535 ;
      RECT 6.815 2.175 6.915 3.135 ;
      RECT 6.215 -48.51 6.565 -48.39 ;
      RECT 6.215 -45.28 6.565 -45.16 ;
      RECT 6.215 -42.05 6.565 -41.93 ;
      RECT 6.215 -38.82 6.565 -38.7 ;
      RECT 6.215 -35.59 6.565 -35.47 ;
      RECT 6.215 -32.36 6.565 -32.24 ;
      RECT 6.215 -29.13 6.565 -29.01 ;
      RECT 6.215 -25.9 6.565 -25.78 ;
      RECT 6.215 -22.67 6.565 -22.55 ;
      RECT 6.215 -19.44 6.565 -19.32 ;
      RECT 6.215 -16.21 6.565 -16.09 ;
      RECT 6.215 -12.98 6.565 -12.86 ;
      RECT 6.215 -9.75 6.565 -9.63 ;
      RECT 6.215 -6.52 6.565 -6.4 ;
      RECT 6.215 -3.29 6.565 -3.17 ;
      RECT 6.215 -0.06 6.565 0.06 ;
      RECT 6.385 -56.495 6.485 -55.535 ;
      RECT 6.385 2.175 6.485 3.135 ;
      RECT 6.28 -59.085 6.45 -58.705 ;
      RECT 6.315 -60.565 6.415 -60.095 ;
      RECT 6.125 -56.495 6.225 -55.535 ;
      RECT 5.875 -56.495 5.975 -55.535 ;
      RECT 5.5 -48.51 5.85 -48.39 ;
      RECT 5.5 -45.28 5.85 -45.16 ;
      RECT 5.5 -42.05 5.85 -41.93 ;
      RECT 5.5 -38.82 5.85 -38.7 ;
      RECT 5.5 -35.59 5.85 -35.47 ;
      RECT 5.5 -32.36 5.85 -32.24 ;
      RECT 5.5 -29.13 5.85 -29.01 ;
      RECT 5.5 -25.9 5.85 -25.78 ;
      RECT 5.5 -22.67 5.85 -22.55 ;
      RECT 5.5 -19.44 5.85 -19.32 ;
      RECT 5.5 -16.21 5.85 -16.09 ;
      RECT 5.5 -12.98 5.85 -12.86 ;
      RECT 5.5 -9.75 5.85 -9.63 ;
      RECT 5.5 -6.52 5.85 -6.4 ;
      RECT 5.5 -3.29 5.85 -3.17 ;
      RECT 5.5 -0.06 5.85 0.06 ;
      RECT 5.615 -56.495 5.715 -55.535 ;
      RECT 5.615 2.175 5.715 3.135 ;
      RECT 5.515 -61.875 5.615 -61.405 ;
      RECT 5.015 -48.51 5.365 -48.39 ;
      RECT 5.015 -45.28 5.365 -45.16 ;
      RECT 5.015 -42.05 5.365 -41.93 ;
      RECT 5.015 -38.82 5.365 -38.7 ;
      RECT 5.015 -35.59 5.365 -35.47 ;
      RECT 5.015 -32.36 5.365 -32.24 ;
      RECT 5.015 -29.13 5.365 -29.01 ;
      RECT 5.015 -25.9 5.365 -25.78 ;
      RECT 5.015 -22.67 5.365 -22.55 ;
      RECT 5.015 -19.44 5.365 -19.32 ;
      RECT 5.015 -16.21 5.365 -16.09 ;
      RECT 5.015 -12.98 5.365 -12.86 ;
      RECT 5.015 -9.75 5.365 -9.63 ;
      RECT 5.015 -6.52 5.365 -6.4 ;
      RECT 5.015 -3.29 5.365 -3.17 ;
      RECT 5.015 -0.06 5.365 0.06 ;
      RECT 5.15 -59.055 5.3 -58.765 ;
      RECT 5.185 -56.495 5.285 -55.535 ;
      RECT 5.185 2.175 5.285 3.135 ;
      RECT 5.165 -60.51 5.265 -59.97 ;
      RECT 4.925 -61.875 5.025 -61.405 ;
      RECT 4.925 -56.495 5.025 -55.535 ;
      RECT 4.675 -53.265 4.775 -52.305 ;
      RECT 4.3 -48.51 4.65 -48.39 ;
      RECT 4.3 -45.28 4.65 -45.16 ;
      RECT 4.3 -42.05 4.65 -41.93 ;
      RECT 4.3 -38.82 4.65 -38.7 ;
      RECT 4.3 -35.59 4.65 -35.47 ;
      RECT 4.3 -32.36 4.65 -32.24 ;
      RECT 4.3 -29.13 4.65 -29.01 ;
      RECT 4.3 -25.9 4.65 -25.78 ;
      RECT 4.3 -22.67 4.65 -22.55 ;
      RECT 4.3 -19.44 4.65 -19.32 ;
      RECT 4.3 -16.21 4.65 -16.09 ;
      RECT 4.3 -12.98 4.65 -12.86 ;
      RECT 4.3 -9.75 4.65 -9.63 ;
      RECT 4.3 -6.52 4.65 -6.4 ;
      RECT 4.3 -3.29 4.65 -3.17 ;
      RECT 4.3 -0.06 4.65 0.06 ;
      RECT 4.415 -53.265 4.515 -52.305 ;
      RECT 4.415 2.175 4.515 3.135 ;
      RECT 4.125 -60.575 4.225 -60.095 ;
      RECT 4.125 -59.085 4.225 -58.615 ;
      RECT 3.815 -48.51 4.165 -48.39 ;
      RECT 3.815 -45.28 4.165 -45.16 ;
      RECT 3.815 -42.05 4.165 -41.93 ;
      RECT 3.815 -38.82 4.165 -38.7 ;
      RECT 3.815 -35.59 4.165 -35.47 ;
      RECT 3.815 -32.36 4.165 -32.24 ;
      RECT 3.815 -29.13 4.165 -29.01 ;
      RECT 3.815 -25.9 4.165 -25.78 ;
      RECT 3.815 -22.67 4.165 -22.55 ;
      RECT 3.815 -19.44 4.165 -19.32 ;
      RECT 3.815 -16.21 4.165 -16.09 ;
      RECT 3.815 -12.98 4.165 -12.86 ;
      RECT 3.815 -9.75 4.165 -9.63 ;
      RECT 3.815 -6.52 4.165 -6.4 ;
      RECT 3.815 -3.29 4.165 -3.17 ;
      RECT 3.815 -0.06 4.165 0.06 ;
      RECT 3.985 -53.265 4.085 -52.305 ;
      RECT 3.985 2.175 4.085 3.135 ;
      RECT 0.085 -56.975 3.865 -56.855 ;
      RECT 3.725 -53.265 3.825 -52.305 ;
      RECT 3.535 -59.07 3.655 -58.69 ;
      RECT 3.535 -60.565 3.635 -60.095 ;
      RECT 3.475 -53.265 3.575 -52.305 ;
      RECT 3.1 -48.51 3.45 -48.39 ;
      RECT 3.1 -45.28 3.45 -45.16 ;
      RECT 3.1 -42.05 3.45 -41.93 ;
      RECT 3.1 -38.82 3.45 -38.7 ;
      RECT 3.1 -35.59 3.45 -35.47 ;
      RECT 3.1 -32.36 3.45 -32.24 ;
      RECT 3.1 -29.13 3.45 -29.01 ;
      RECT 3.1 -25.9 3.45 -25.78 ;
      RECT 3.1 -22.67 3.45 -22.55 ;
      RECT 3.1 -19.44 3.45 -19.32 ;
      RECT 3.1 -16.21 3.45 -16.09 ;
      RECT 3.1 -12.98 3.45 -12.86 ;
      RECT 3.1 -9.75 3.45 -9.63 ;
      RECT 3.1 -6.52 3.45 -6.4 ;
      RECT 3.1 -3.29 3.45 -3.17 ;
      RECT 3.1 -0.06 3.45 0.06 ;
      RECT 3.215 -53.265 3.315 -52.305 ;
      RECT 3.215 2.175 3.315 3.135 ;
      RECT 2.945 -57.915 3.08 -57.595 ;
      RECT 2.615 -48.51 2.965 -48.39 ;
      RECT 2.615 -45.28 2.965 -45.16 ;
      RECT 2.615 -42.05 2.965 -41.93 ;
      RECT 2.615 -38.82 2.965 -38.7 ;
      RECT 2.615 -35.59 2.965 -35.47 ;
      RECT 2.615 -32.36 2.965 -32.24 ;
      RECT 2.615 -29.13 2.965 -29.01 ;
      RECT 2.615 -25.9 2.965 -25.78 ;
      RECT 2.615 -22.67 2.965 -22.55 ;
      RECT 2.615 -19.44 2.965 -19.32 ;
      RECT 2.615 -16.21 2.965 -16.09 ;
      RECT 2.615 -12.98 2.965 -12.86 ;
      RECT 2.615 -9.75 2.965 -9.63 ;
      RECT 2.615 -6.52 2.965 -6.4 ;
      RECT 2.615 -3.29 2.965 -3.17 ;
      RECT 2.615 -0.06 2.965 0.06 ;
      RECT 2.785 -53.265 2.885 -52.305 ;
      RECT 2.785 2.175 2.885 3.135 ;
      RECT 2.61 -57.915 2.755 -57.595 ;
      RECT 2.525 -53.265 2.625 -52.305 ;
      RECT 2.275 -56.495 2.375 -55.535 ;
      RECT 1.9 -48.51 2.25 -48.39 ;
      RECT 1.9 -45.28 2.25 -45.16 ;
      RECT 1.9 -42.05 2.25 -41.93 ;
      RECT 1.9 -38.82 2.25 -38.7 ;
      RECT 1.9 -35.59 2.25 -35.47 ;
      RECT 1.9 -32.36 2.25 -32.24 ;
      RECT 1.9 -29.13 2.25 -29.01 ;
      RECT 1.9 -25.9 2.25 -25.78 ;
      RECT 1.9 -22.67 2.25 -22.55 ;
      RECT 1.9 -19.44 2.25 -19.32 ;
      RECT 1.9 -16.21 2.25 -16.09 ;
      RECT 1.9 -12.98 2.25 -12.86 ;
      RECT 1.9 -9.75 2.25 -9.63 ;
      RECT 1.9 -6.52 2.25 -6.4 ;
      RECT 1.9 -3.29 2.25 -3.17 ;
      RECT 1.9 -0.06 2.25 0.06 ;
      RECT 2.105 -60.575 2.205 -60.095 ;
      RECT 2.105 -59.085 2.205 -58.615 ;
      RECT 2.015 -56.495 2.115 -55.535 ;
      RECT 2.015 2.175 2.115 3.135 ;
      RECT 1.415 -48.51 1.765 -48.39 ;
      RECT 1.415 -45.28 1.765 -45.16 ;
      RECT 1.415 -42.05 1.765 -41.93 ;
      RECT 1.415 -38.82 1.765 -38.7 ;
      RECT 1.415 -35.59 1.765 -35.47 ;
      RECT 1.415 -32.36 1.765 -32.24 ;
      RECT 1.415 -29.13 1.765 -29.01 ;
      RECT 1.415 -25.9 1.765 -25.78 ;
      RECT 1.415 -22.67 1.765 -22.55 ;
      RECT 1.415 -19.44 1.765 -19.32 ;
      RECT 1.415 -16.21 1.765 -16.09 ;
      RECT 1.415 -12.98 1.765 -12.86 ;
      RECT 1.415 -9.75 1.765 -9.63 ;
      RECT 1.415 -6.52 1.765 -6.4 ;
      RECT 1.415 -3.29 1.765 -3.17 ;
      RECT 1.415 -0.06 1.765 0.06 ;
      RECT 1.585 -56.495 1.685 -55.535 ;
      RECT 1.585 2.175 1.685 3.135 ;
      RECT 1.48 -59.085 1.65 -58.705 ;
      RECT 1.515 -60.565 1.615 -60.095 ;
      RECT 1.325 -56.495 1.425 -55.535 ;
      RECT 1.075 -56.495 1.175 -55.535 ;
      RECT 0.7 -48.51 1.05 -48.39 ;
      RECT 0.7 -45.28 1.05 -45.16 ;
      RECT 0.7 -42.05 1.05 -41.93 ;
      RECT 0.7 -38.82 1.05 -38.7 ;
      RECT 0.7 -35.59 1.05 -35.47 ;
      RECT 0.7 -32.36 1.05 -32.24 ;
      RECT 0.7 -29.13 1.05 -29.01 ;
      RECT 0.7 -25.9 1.05 -25.78 ;
      RECT 0.7 -22.67 1.05 -22.55 ;
      RECT 0.7 -19.44 1.05 -19.32 ;
      RECT 0.7 -16.21 1.05 -16.09 ;
      RECT 0.7 -12.98 1.05 -12.86 ;
      RECT 0.7 -9.75 1.05 -9.63 ;
      RECT 0.7 -6.52 1.05 -6.4 ;
      RECT 0.7 -3.29 1.05 -3.17 ;
      RECT 0.7 -0.06 1.05 0.06 ;
      RECT 0.815 -56.495 0.915 -55.535 ;
      RECT 0.815 2.175 0.915 3.135 ;
      RECT 0.715 -61.875 0.815 -61.405 ;
      RECT 0.215 -48.51 0.565 -48.39 ;
      RECT 0.215 -45.28 0.565 -45.16 ;
      RECT 0.215 -42.05 0.565 -41.93 ;
      RECT 0.215 -38.82 0.565 -38.7 ;
      RECT 0.215 -35.59 0.565 -35.47 ;
      RECT 0.215 -32.36 0.565 -32.24 ;
      RECT 0.215 -29.13 0.565 -29.01 ;
      RECT 0.215 -25.9 0.565 -25.78 ;
      RECT 0.215 -22.67 0.565 -22.55 ;
      RECT 0.215 -19.44 0.565 -19.32 ;
      RECT 0.215 -16.21 0.565 -16.09 ;
      RECT 0.215 -12.98 0.565 -12.86 ;
      RECT 0.215 -9.75 0.565 -9.63 ;
      RECT 0.215 -6.52 0.565 -6.4 ;
      RECT 0.215 -3.29 0.565 -3.17 ;
      RECT 0.215 -0.06 0.565 0.06 ;
      RECT 0.35 -59.055 0.5 -58.765 ;
      RECT 0.385 -56.495 0.485 -55.535 ;
      RECT 0.385 2.175 0.485 3.135 ;
      RECT 0.365 -60.51 0.465 -59.97 ;
      RECT 0.125 -61.875 0.225 -61.405 ;
      RECT 0.125 -56.495 0.225 -55.535 ;
      RECT -0.765 -55.975 -0.665 -55.555 ;
      RECT -0.765 -51.215 -0.665 -50.615 ;
      RECT -0.765 -49.515 -0.665 -48.915 ;
      RECT -0.765 -44.575 -0.665 -44.155 ;
      RECT -0.765 -43.055 -0.665 -42.635 ;
      RECT -0.765 -38.295 -0.665 -37.695 ;
      RECT -0.765 -36.595 -0.665 -35.995 ;
      RECT -0.765 -31.655 -0.665 -31.235 ;
      RECT -0.765 -30.135 -0.665 -29.715 ;
      RECT -0.765 -25.375 -0.665 -24.775 ;
      RECT -0.765 -23.675 -0.665 -23.075 ;
      RECT -0.765 -18.735 -0.665 -18.315 ;
      RECT -0.765 -17.215 -0.665 -16.795 ;
      RECT -0.765 -12.455 -0.665 -11.855 ;
      RECT -0.765 -10.755 -0.665 -10.155 ;
      RECT -0.765 -5.815 -0.665 -5.395 ;
      RECT -0.765 -4.295 -0.665 -3.875 ;
      RECT -0.765 0.465 -0.665 1.065 ;
      RECT -1.845 -51.73 -0.76 -51.63 ;
      RECT -1.845 -48.5 -0.76 -48.4 ;
      RECT -1.845 -38.81 -0.76 -38.71 ;
      RECT -1.845 -35.58 -0.76 -35.48 ;
      RECT -1.845 -25.89 -0.76 -25.79 ;
      RECT -1.845 -22.66 -0.76 -22.56 ;
      RECT -1.845 -12.97 -0.76 -12.87 ;
      RECT -1.845 -9.74 -0.76 -9.64 ;
      RECT -1.845 -0.05 -0.76 0.05 ;
      RECT -1.285 -55.975 -1.185 -55.375 ;
      RECT -1.285 -51.215 -1.185 -50.615 ;
      RECT -1.285 -49.515 -1.185 -48.915 ;
      RECT -1.285 -44.755 -1.185 -44.155 ;
      RECT -1.285 -43.055 -1.185 -42.455 ;
      RECT -1.285 -38.295 -1.185 -37.695 ;
      RECT -1.285 -36.595 -1.185 -35.995 ;
      RECT -1.285 -31.835 -1.185 -31.235 ;
      RECT -1.285 -30.135 -1.185 -29.535 ;
      RECT -1.285 -25.375 -1.185 -24.775 ;
      RECT -1.285 -23.675 -1.185 -23.075 ;
      RECT -1.285 -18.915 -1.185 -18.315 ;
      RECT -1.285 -17.215 -1.185 -16.615 ;
      RECT -1.285 -12.455 -1.185 -11.855 ;
      RECT -1.285 -10.755 -1.185 -10.155 ;
      RECT -1.285 -5.995 -1.185 -5.395 ;
      RECT -1.285 -4.295 -1.185 -3.695 ;
      RECT -1.285 0.465 -1.185 1.065 ;
      RECT -8.605 -52.975 -1.28 -52.875 ;
      RECT -16.405 -46.375 -1.28 -46.275 ;
      RECT -16.405 -40.935 -1.28 -40.835 ;
      RECT -16.405 -33.455 -1.28 -33.355 ;
      RECT -16.405 -28.015 -1.28 -27.915 ;
      RECT -16.405 -20.535 -1.28 -20.435 ;
      RECT -16.405 -15.095 -1.28 -14.995 ;
      RECT -16.405 -7.615 -1.28 -7.515 ;
      RECT -16.405 -2.175 -1.28 -2.075 ;
      RECT -1.545 -55.975 -1.445 -55.375 ;
      RECT -1.545 -44.755 -1.445 -44.155 ;
      RECT -1.545 -43.055 -1.445 -42.455 ;
      RECT -1.545 -31.835 -1.445 -31.235 ;
      RECT -1.545 -30.135 -1.445 -29.535 ;
      RECT -1.545 -18.915 -1.445 -18.315 ;
      RECT -1.545 -17.215 -1.445 -16.615 ;
      RECT -1.545 -5.995 -1.445 -5.395 ;
      RECT -1.545 -4.295 -1.445 -3.695 ;
      RECT -5.905 -52.315 -1.54 -52.215 ;
      RECT -5.905 -47.695 -1.54 -47.595 ;
      RECT -5.905 -39.615 -1.54 -39.515 ;
      RECT -5.905 -34.775 -1.54 -34.675 ;
      RECT -5.905 -26.695 -1.54 -26.595 ;
      RECT -5.905 -21.855 -1.54 -21.755 ;
      RECT -5.905 -13.775 -1.54 -13.675 ;
      RECT -5.905 -8.935 -1.54 -8.835 ;
      RECT -5.905 -0.855 -1.54 -0.755 ;
      RECT -1.805 -51.215 -1.705 -50.615 ;
      RECT -1.805 -49.515 -1.705 -48.915 ;
      RECT -1.805 -38.295 -1.705 -37.695 ;
      RECT -1.805 -36.595 -1.705 -35.995 ;
      RECT -1.805 -25.375 -1.705 -24.775 ;
      RECT -1.805 -23.675 -1.705 -23.075 ;
      RECT -1.805 -12.455 -1.705 -11.855 ;
      RECT -1.805 -10.755 -1.705 -10.155 ;
      RECT -1.805 0.465 -1.705 1.065 ;
      RECT -2.065 -55.975 -1.965 -55.555 ;
      RECT -2.065 -51.215 -1.965 -50.615 ;
      RECT -2.065 -49.515 -1.965 -48.915 ;
      RECT -2.065 -44.575 -1.965 -44.155 ;
      RECT -2.065 -43.055 -1.965 -42.635 ;
      RECT -2.065 -38.295 -1.965 -37.695 ;
      RECT -2.065 -36.595 -1.965 -35.995 ;
      RECT -2.065 -31.655 -1.965 -31.235 ;
      RECT -2.065 -30.135 -1.965 -29.715 ;
      RECT -2.065 -25.375 -1.965 -24.775 ;
      RECT -2.065 -23.675 -1.965 -23.075 ;
      RECT -2.065 -18.735 -1.965 -18.315 ;
      RECT -2.065 -17.215 -1.965 -16.795 ;
      RECT -2.065 -12.455 -1.965 -11.855 ;
      RECT -2.065 -10.755 -1.965 -10.155 ;
      RECT -2.065 -5.815 -1.965 -5.395 ;
      RECT -2.065 -4.295 -1.965 -3.875 ;
      RECT -2.065 0.465 -1.965 1.065 ;
      RECT -3.145 -51.73 -2.06 -51.63 ;
      RECT -3.145 -48.5 -2.06 -48.4 ;
      RECT -3.145 -38.81 -2.06 -38.71 ;
      RECT -3.145 -35.58 -2.06 -35.48 ;
      RECT -3.145 -25.89 -2.06 -25.79 ;
      RECT -3.145 -22.66 -2.06 -22.56 ;
      RECT -3.145 -12.97 -2.06 -12.87 ;
      RECT -3.145 -9.74 -2.06 -9.64 ;
      RECT -3.145 -0.05 -2.06 0.05 ;
      RECT -2.585 -55.975 -2.485 -55.375 ;
      RECT -2.585 -51.215 -2.485 -50.615 ;
      RECT -2.585 -49.515 -2.485 -48.915 ;
      RECT -2.585 -44.755 -2.485 -44.155 ;
      RECT -2.585 -43.055 -2.485 -42.455 ;
      RECT -2.585 -38.295 -2.485 -37.695 ;
      RECT -2.585 -36.595 -2.485 -35.995 ;
      RECT -2.585 -31.835 -2.485 -31.235 ;
      RECT -2.585 -30.135 -2.485 -29.535 ;
      RECT -2.585 -25.375 -2.485 -24.775 ;
      RECT -2.585 -23.675 -2.485 -23.075 ;
      RECT -2.585 -18.915 -2.485 -18.315 ;
      RECT -2.585 -17.215 -2.485 -16.615 ;
      RECT -2.585 -12.455 -2.485 -11.855 ;
      RECT -2.585 -10.755 -2.485 -10.155 ;
      RECT -2.585 -5.995 -2.485 -5.395 ;
      RECT -2.585 -4.295 -2.485 -3.695 ;
      RECT -2.585 0.465 -2.485 1.065 ;
      RECT -9.905 -52.755 -2.58 -52.655 ;
      RECT -21.605 -46.595 -2.58 -46.495 ;
      RECT -21.605 -40.715 -2.58 -40.615 ;
      RECT -21.605 -33.675 -2.58 -33.575 ;
      RECT -21.605 -27.795 -2.58 -27.695 ;
      RECT -21.605 -20.755 -2.58 -20.655 ;
      RECT -21.605 -14.875 -2.58 -14.775 ;
      RECT -21.605 -7.835 -2.58 -7.735 ;
      RECT -21.605 -1.955 -2.58 -1.855 ;
      RECT -2.845 -55.975 -2.745 -55.375 ;
      RECT -2.845 -44.755 -2.745 -44.155 ;
      RECT -2.845 -43.055 -2.745 -42.455 ;
      RECT -2.845 -31.835 -2.745 -31.235 ;
      RECT -2.845 -30.135 -2.745 -29.535 ;
      RECT -2.845 -18.915 -2.745 -18.315 ;
      RECT -2.845 -17.215 -2.745 -16.615 ;
      RECT -2.845 -5.995 -2.745 -5.395 ;
      RECT -2.845 -4.295 -2.745 -3.695 ;
      RECT -3.105 -51.215 -3.005 -50.615 ;
      RECT -3.105 -49.515 -3.005 -48.915 ;
      RECT -3.105 -38.295 -3.005 -37.695 ;
      RECT -3.105 -36.595 -3.005 -35.995 ;
      RECT -3.105 -25.375 -3.005 -24.775 ;
      RECT -3.105 -23.675 -3.005 -23.075 ;
      RECT -3.105 -12.455 -3.005 -11.855 ;
      RECT -3.105 -10.755 -3.005 -10.155 ;
      RECT -3.105 0.465 -3.005 1.065 ;
      RECT -3.365 -55.975 -3.265 -55.555 ;
      RECT -3.365 -51.215 -3.265 -50.615 ;
      RECT -3.365 -49.515 -3.265 -48.915 ;
      RECT -3.365 -44.575 -3.265 -44.155 ;
      RECT -3.365 -43.055 -3.265 -42.635 ;
      RECT -3.365 -38.295 -3.265 -37.695 ;
      RECT -3.365 -36.595 -3.265 -35.995 ;
      RECT -3.365 -31.655 -3.265 -31.235 ;
      RECT -3.365 -30.135 -3.265 -29.715 ;
      RECT -3.365 -25.375 -3.265 -24.775 ;
      RECT -3.365 -23.675 -3.265 -23.075 ;
      RECT -3.365 -18.735 -3.265 -18.315 ;
      RECT -3.365 -17.215 -3.265 -16.795 ;
      RECT -3.365 -12.455 -3.265 -11.855 ;
      RECT -3.365 -10.755 -3.265 -10.155 ;
      RECT -3.365 -5.815 -3.265 -5.395 ;
      RECT -3.365 -4.295 -3.265 -3.875 ;
      RECT -3.365 0.465 -3.265 1.065 ;
      RECT -4.445 -51.73 -3.36 -51.63 ;
      RECT -4.445 -48.5 -3.36 -48.4 ;
      RECT -4.445 -38.81 -3.36 -38.71 ;
      RECT -4.445 -35.58 -3.36 -35.48 ;
      RECT -4.445 -25.89 -3.36 -25.79 ;
      RECT -4.445 -22.66 -3.36 -22.56 ;
      RECT -4.445 -12.97 -3.36 -12.87 ;
      RECT -4.445 -9.74 -3.36 -9.64 ;
      RECT -4.445 -0.05 -3.36 0.05 ;
      RECT -3.885 -55.975 -3.785 -55.375 ;
      RECT -3.885 -51.215 -3.785 -50.615 ;
      RECT -3.885 -49.515 -3.785 -48.915 ;
      RECT -3.885 -44.755 -3.785 -44.155 ;
      RECT -3.885 -43.055 -3.785 -42.455 ;
      RECT -3.885 -38.295 -3.785 -37.695 ;
      RECT -3.885 -36.595 -3.785 -35.995 ;
      RECT -3.885 -31.835 -3.785 -31.235 ;
      RECT -3.885 -30.135 -3.785 -29.535 ;
      RECT -3.885 -25.375 -3.785 -24.775 ;
      RECT -3.885 -23.675 -3.785 -23.075 ;
      RECT -3.885 -18.915 -3.785 -18.315 ;
      RECT -3.885 -17.215 -3.785 -16.615 ;
      RECT -3.885 -12.455 -3.785 -11.855 ;
      RECT -3.885 -10.755 -3.785 -10.155 ;
      RECT -3.885 -5.995 -3.785 -5.395 ;
      RECT -3.885 -4.295 -3.785 -3.695 ;
      RECT -3.885 0.465 -3.785 1.065 ;
      RECT -6.005 -52.535 -3.88 -52.435 ;
      RECT -6.005 -46.815 -3.88 -46.715 ;
      RECT -6.005 -40.495 -3.88 -40.395 ;
      RECT -6.005 -33.895 -3.88 -33.795 ;
      RECT -6.005 -27.575 -3.88 -27.475 ;
      RECT -6.005 -20.975 -3.88 -20.875 ;
      RECT -6.005 -14.655 -3.88 -14.555 ;
      RECT -6.005 -8.055 -3.88 -7.955 ;
      RECT -6.005 -1.735 -3.88 -1.635 ;
      RECT -4.145 -55.975 -4.045 -55.375 ;
      RECT -4.145 -44.755 -4.045 -44.155 ;
      RECT -4.145 -43.055 -4.045 -42.455 ;
      RECT -4.145 -31.835 -4.045 -31.235 ;
      RECT -4.145 -30.135 -4.045 -29.535 ;
      RECT -4.145 -18.915 -4.045 -18.315 ;
      RECT -4.145 -17.215 -4.045 -16.615 ;
      RECT -4.145 -5.995 -4.045 -5.395 ;
      RECT -4.145 -4.295 -4.045 -3.695 ;
      RECT -4.405 -51.215 -4.305 -50.615 ;
      RECT -4.405 -49.515 -4.305 -48.915 ;
      RECT -4.405 -38.295 -4.305 -37.695 ;
      RECT -4.405 -36.595 -4.305 -35.995 ;
      RECT -4.405 -25.375 -4.305 -24.775 ;
      RECT -4.405 -23.675 -4.305 -23.075 ;
      RECT -4.405 -12.455 -4.305 -11.855 ;
      RECT -4.405 -10.755 -4.305 -10.155 ;
      RECT -4.405 0.465 -4.305 1.065 ;
      RECT -4.665 -55.975 -4.565 -55.555 ;
      RECT -4.665 -51.215 -4.565 -50.615 ;
      RECT -4.665 -49.515 -4.565 -48.915 ;
      RECT -4.665 -44.575 -4.565 -44.155 ;
      RECT -4.665 -43.055 -4.565 -42.635 ;
      RECT -4.665 -38.295 -4.565 -37.695 ;
      RECT -4.665 -36.595 -4.565 -35.995 ;
      RECT -4.665 -31.655 -4.565 -31.235 ;
      RECT -4.665 -30.135 -4.565 -29.715 ;
      RECT -4.665 -25.375 -4.565 -24.775 ;
      RECT -4.665 -23.675 -4.565 -23.075 ;
      RECT -4.665 -18.735 -4.565 -18.315 ;
      RECT -4.665 -17.215 -4.565 -16.795 ;
      RECT -4.665 -12.455 -4.565 -11.855 ;
      RECT -4.665 -10.755 -4.565 -10.155 ;
      RECT -4.665 -5.815 -4.565 -5.395 ;
      RECT -4.665 -4.295 -4.565 -3.875 ;
      RECT -4.665 0.465 -4.565 1.065 ;
      RECT -5.745 -51.73 -4.66 -51.63 ;
      RECT -5.745 -48.5 -4.66 -48.4 ;
      RECT -5.745 -38.81 -4.66 -38.71 ;
      RECT -5.745 -35.58 -4.66 -35.48 ;
      RECT -5.745 -25.89 -4.66 -25.79 ;
      RECT -5.745 -22.66 -4.66 -22.56 ;
      RECT -5.745 -12.97 -4.66 -12.87 ;
      RECT -5.745 -9.74 -4.66 -9.64 ;
      RECT -5.745 -0.05 -4.66 0.05 ;
      RECT -5.185 -55.975 -5.085 -55.375 ;
      RECT -5.185 -51.215 -5.085 -50.615 ;
      RECT -5.185 -49.515 -5.085 -48.915 ;
      RECT -5.185 -44.755 -5.085 -44.155 ;
      RECT -5.185 -43.055 -5.085 -42.455 ;
      RECT -5.185 -38.295 -5.085 -37.695 ;
      RECT -5.185 -36.595 -5.085 -35.995 ;
      RECT -5.185 -31.835 -5.085 -31.235 ;
      RECT -5.185 -30.135 -5.085 -29.535 ;
      RECT -5.185 -25.375 -5.085 -24.775 ;
      RECT -5.185 -23.675 -5.085 -23.075 ;
      RECT -5.185 -18.915 -5.085 -18.315 ;
      RECT -5.185 -17.215 -5.085 -16.615 ;
      RECT -5.185 -12.455 -5.085 -11.855 ;
      RECT -5.185 -10.755 -5.085 -10.155 ;
      RECT -5.185 -5.995 -5.085 -5.395 ;
      RECT -5.185 -4.295 -5.085 -3.695 ;
      RECT -5.185 0.465 -5.085 1.065 ;
      RECT -7.305 -52.095 -5.18 -51.995 ;
      RECT -11.205 -48.135 -5.18 -48.035 ;
      RECT -11.205 -39.175 -5.18 -39.075 ;
      RECT -11.205 -35.215 -5.18 -35.115 ;
      RECT -11.205 -26.255 -5.18 -26.155 ;
      RECT -11.205 -22.295 -5.18 -22.195 ;
      RECT -11.205 -13.335 -5.18 -13.235 ;
      RECT -11.205 -9.375 -5.18 -9.275 ;
      RECT -11.205 -0.415 -5.18 -0.315 ;
      RECT -5.445 -55.975 -5.345 -55.375 ;
      RECT -5.445 -44.755 -5.345 -44.155 ;
      RECT -5.445 -43.055 -5.345 -42.455 ;
      RECT -5.445 -31.835 -5.345 -31.235 ;
      RECT -5.445 -30.135 -5.345 -29.535 ;
      RECT -5.445 -18.915 -5.345 -18.315 ;
      RECT -5.445 -17.215 -5.345 -16.615 ;
      RECT -5.445 -5.995 -5.345 -5.395 ;
      RECT -5.445 -4.295 -5.345 -3.695 ;
      RECT -5.705 -51.215 -5.605 -50.615 ;
      RECT -5.705 -49.515 -5.605 -48.915 ;
      RECT -5.705 -38.295 -5.605 -37.695 ;
      RECT -5.705 -36.595 -5.605 -35.995 ;
      RECT -5.705 -25.375 -5.605 -24.775 ;
      RECT -5.705 -23.675 -5.605 -23.075 ;
      RECT -5.705 -12.455 -5.605 -11.855 ;
      RECT -5.705 -10.755 -5.605 -10.155 ;
      RECT -5.705 0.465 -5.605 1.065 ;
      RECT -5.965 -55.975 -5.865 -55.555 ;
      RECT -5.965 -51.215 -5.865 -50.615 ;
      RECT -5.965 -49.515 -5.865 -48.915 ;
      RECT -5.965 -44.575 -5.865 -44.155 ;
      RECT -5.965 -43.055 -5.865 -42.635 ;
      RECT -5.965 -38.295 -5.865 -37.695 ;
      RECT -5.965 -36.595 -5.865 -35.995 ;
      RECT -5.965 -31.655 -5.865 -31.235 ;
      RECT -5.965 -30.135 -5.865 -29.715 ;
      RECT -5.965 -25.375 -5.865 -24.775 ;
      RECT -5.965 -23.675 -5.865 -23.075 ;
      RECT -5.965 -18.735 -5.865 -18.315 ;
      RECT -5.965 -17.215 -5.865 -16.795 ;
      RECT -5.965 -12.455 -5.865 -11.855 ;
      RECT -5.965 -10.755 -5.865 -10.155 ;
      RECT -5.965 -5.815 -5.865 -5.395 ;
      RECT -5.965 -4.295 -5.865 -3.875 ;
      RECT -5.965 0.465 -5.865 1.065 ;
      RECT -6.485 -55.975 -6.385 -55.375 ;
      RECT -6.485 -44.755 -6.385 -44.155 ;
      RECT -6.485 -43.055 -6.385 -42.455 ;
      RECT -6.485 -31.835 -6.385 -31.235 ;
      RECT -6.485 -30.135 -6.385 -29.535 ;
      RECT -6.485 -18.915 -6.385 -18.315 ;
      RECT -6.485 -17.215 -6.385 -16.615 ;
      RECT -6.485 -5.995 -6.385 -5.395 ;
      RECT -6.485 -4.295 -6.385 -3.695 ;
      RECT -7.305 -47.035 -6.48 -46.935 ;
      RECT -7.305 -40.275 -6.48 -40.175 ;
      RECT -7.305 -34.115 -6.48 -34.015 ;
      RECT -7.305 -27.355 -6.48 -27.255 ;
      RECT -7.305 -21.195 -6.48 -21.095 ;
      RECT -7.305 -14.435 -6.48 -14.335 ;
      RECT -7.305 -8.275 -6.48 -8.175 ;
      RECT -7.305 -1.515 -6.48 -1.415 ;
      RECT -6.745 -55.975 -6.645 -55.375 ;
      RECT -6.745 -44.755 -6.645 -44.155 ;
      RECT -6.745 -43.055 -6.645 -42.455 ;
      RECT -6.745 -31.835 -6.645 -31.235 ;
      RECT -6.745 -30.135 -6.645 -29.535 ;
      RECT -6.745 -18.915 -6.645 -18.315 ;
      RECT -6.745 -17.215 -6.645 -16.615 ;
      RECT -6.745 -5.995 -6.645 -5.395 ;
      RECT -6.745 -4.295 -6.645 -3.695 ;
      RECT -29.865 -21.415 -6.74 -21.315 ;
      RECT -29.865 -14.215 -6.74 -14.115 ;
      RECT -29.865 -8.495 -6.74 -8.395 ;
      RECT -29.865 -1.295 -6.74 -1.195 ;
      RECT -7.265 -55.975 -7.165 -55.555 ;
      RECT -7.265 -51.215 -7.165 -50.615 ;
      RECT -7.265 -49.515 -7.165 -48.915 ;
      RECT -7.265 -44.575 -7.165 -44.155 ;
      RECT -7.265 -43.055 -7.165 -42.635 ;
      RECT -7.265 -38.295 -7.165 -37.695 ;
      RECT -7.265 -36.595 -7.165 -35.995 ;
      RECT -7.265 -31.655 -7.165 -31.235 ;
      RECT -7.265 -30.135 -7.165 -29.715 ;
      RECT -7.265 -25.375 -7.165 -24.775 ;
      RECT -7.265 -23.675 -7.165 -23.075 ;
      RECT -7.265 -18.735 -7.165 -18.315 ;
      RECT -7.265 -17.215 -7.165 -16.795 ;
      RECT -7.265 -12.455 -7.165 -11.855 ;
      RECT -7.265 -10.755 -7.165 -10.155 ;
      RECT -7.265 -5.815 -7.165 -5.395 ;
      RECT -7.265 -4.295 -7.165 -3.875 ;
      RECT -7.265 0.465 -7.165 1.065 ;
      RECT -7.785 -55.975 -7.685 -55.375 ;
      RECT -7.785 -44.755 -7.685 -44.155 ;
      RECT -7.785 -43.055 -7.685 -42.455 ;
      RECT -7.785 -31.835 -7.685 -31.235 ;
      RECT -7.785 -30.135 -7.685 -29.535 ;
      RECT -7.785 -18.915 -7.685 -18.315 ;
      RECT -7.785 -17.215 -7.685 -16.615 ;
      RECT -7.785 -5.995 -7.685 -5.395 ;
      RECT -7.785 -4.295 -7.685 -3.695 ;
      RECT -8.605 -46.815 -7.78 -46.715 ;
      RECT -8.605 -40.495 -7.78 -40.395 ;
      RECT -8.605 -33.895 -7.78 -33.795 ;
      RECT -8.605 -27.575 -7.78 -27.475 ;
      RECT -8.605 -20.975 -7.78 -20.875 ;
      RECT -8.605 -14.655 -7.78 -14.555 ;
      RECT -8.605 -8.055 -7.78 -7.955 ;
      RECT -8.605 -1.735 -7.78 -1.635 ;
      RECT -8.045 -55.975 -7.945 -55.375 ;
      RECT -8.045 -44.755 -7.945 -44.155 ;
      RECT -8.045 -43.055 -7.945 -42.455 ;
      RECT -8.045 -31.835 -7.945 -31.235 ;
      RECT -8.045 -30.135 -7.945 -29.535 ;
      RECT -8.045 -18.915 -7.945 -18.315 ;
      RECT -8.045 -17.215 -7.945 -16.615 ;
      RECT -8.045 -5.995 -7.945 -5.395 ;
      RECT -8.045 -4.295 -7.945 -3.695 ;
      RECT -12.465 -51.655 -8.04 -51.555 ;
      RECT -9.905 -47.035 -8.04 -46.935 ;
      RECT -9.905 -40.275 -8.04 -40.175 ;
      RECT -9.905 -34.115 -8.04 -34.015 ;
      RECT -9.905 -27.355 -8.04 -27.255 ;
      RECT -9.905 -21.195 -8.04 -21.095 ;
      RECT -9.905 -14.435 -8.04 -14.335 ;
      RECT -9.905 -8.275 -8.04 -8.175 ;
      RECT -9.905 -1.515 -8.04 -1.415 ;
      RECT -8.565 -55.975 -8.465 -55.555 ;
      RECT -8.565 -51.215 -8.465 -50.615 ;
      RECT -8.565 -49.515 -8.465 -48.915 ;
      RECT -8.565 -44.575 -8.465 -44.155 ;
      RECT -8.565 -43.055 -8.465 -42.635 ;
      RECT -8.565 -38.295 -8.465 -37.695 ;
      RECT -8.565 -36.595 -8.465 -35.995 ;
      RECT -8.565 -31.655 -8.465 -31.235 ;
      RECT -8.565 -30.135 -8.465 -29.715 ;
      RECT -8.565 -25.375 -8.465 -24.775 ;
      RECT -8.565 -23.675 -8.465 -23.075 ;
      RECT -8.565 -18.735 -8.465 -18.315 ;
      RECT -8.565 -17.215 -8.465 -16.795 ;
      RECT -8.565 -12.455 -8.465 -11.855 ;
      RECT -8.565 -10.755 -8.465 -10.155 ;
      RECT -8.565 -5.815 -8.465 -5.395 ;
      RECT -8.565 -4.295 -8.465 -3.875 ;
      RECT -8.565 0.465 -8.465 1.065 ;
      RECT -9.085 -55.975 -8.985 -55.375 ;
      RECT -9.085 -44.755 -8.985 -44.155 ;
      RECT -9.085 -43.055 -8.985 -42.455 ;
      RECT -9.085 -31.835 -8.985 -31.235 ;
      RECT -9.085 -30.135 -8.985 -29.535 ;
      RECT -9.085 -18.915 -8.985 -18.315 ;
      RECT -9.085 -17.215 -8.985 -16.615 ;
      RECT -9.085 -5.995 -8.985 -5.395 ;
      RECT -9.085 -4.295 -8.985 -3.695 ;
      RECT -12.465 -52.095 -9.08 -51.995 ;
      RECT -29.865 -34.555 -9.08 -34.455 ;
      RECT -29.865 -26.915 -9.08 -26.815 ;
      RECT -29.865 -8.715 -9.08 -8.615 ;
      RECT -29.865 -1.075 -9.08 -0.975 ;
      RECT -9.345 -55.975 -9.245 -55.375 ;
      RECT -9.345 -44.755 -9.245 -44.155 ;
      RECT -9.345 -43.055 -9.245 -42.455 ;
      RECT -9.345 -31.835 -9.245 -31.235 ;
      RECT -9.345 -30.135 -9.245 -29.535 ;
      RECT -9.345 -18.915 -9.245 -18.315 ;
      RECT -9.345 -17.215 -9.245 -16.615 ;
      RECT -9.345 -5.995 -9.245 -5.395 ;
      RECT -9.345 -4.295 -9.245 -3.695 ;
      RECT -29.865 -39.615 -9.34 -39.515 ;
      RECT -29.865 -26.695 -9.34 -26.595 ;
      RECT -29.865 -13.775 -9.34 -13.675 ;
      RECT -29.865 -0.855 -9.34 -0.755 ;
      RECT -9.865 -55.975 -9.765 -55.555 ;
      RECT -9.865 -51.215 -9.765 -50.615 ;
      RECT -9.865 -49.515 -9.765 -48.915 ;
      RECT -9.865 -44.575 -9.765 -44.155 ;
      RECT -9.865 -43.055 -9.765 -42.635 ;
      RECT -9.865 -38.295 -9.765 -37.695 ;
      RECT -9.865 -36.595 -9.765 -35.995 ;
      RECT -9.865 -31.655 -9.765 -31.235 ;
      RECT -9.865 -30.135 -9.765 -29.715 ;
      RECT -9.865 -25.375 -9.765 -24.775 ;
      RECT -9.865 -23.675 -9.765 -23.075 ;
      RECT -9.865 -18.735 -9.765 -18.315 ;
      RECT -9.865 -17.215 -9.765 -16.795 ;
      RECT -9.865 -12.455 -9.765 -11.855 ;
      RECT -9.865 -10.755 -9.765 -10.155 ;
      RECT -9.865 -5.815 -9.765 -5.395 ;
      RECT -9.865 -4.295 -9.765 -3.875 ;
      RECT -9.865 0.465 -9.765 1.065 ;
      RECT -10.385 -55.975 -10.285 -55.375 ;
      RECT -10.385 -44.755 -10.285 -44.155 ;
      RECT -10.385 -43.055 -10.285 -42.455 ;
      RECT -10.385 -31.835 -10.285 -31.235 ;
      RECT -10.385 -30.135 -10.285 -29.535 ;
      RECT -10.385 -18.915 -10.285 -18.315 ;
      RECT -10.385 -17.215 -10.285 -16.615 ;
      RECT -10.385 -5.995 -10.285 -5.395 ;
      RECT -10.385 -4.295 -10.285 -3.695 ;
      RECT -10.645 -55.975 -10.545 -55.375 ;
      RECT -10.645 -44.755 -10.545 -44.155 ;
      RECT -10.645 -43.055 -10.545 -42.455 ;
      RECT -10.645 -31.835 -10.545 -31.235 ;
      RECT -10.645 -30.135 -10.545 -29.535 ;
      RECT -10.645 -18.915 -10.545 -18.315 ;
      RECT -10.645 -17.215 -10.545 -16.615 ;
      RECT -10.645 -5.995 -10.545 -5.395 ;
      RECT -10.645 -4.295 -10.545 -3.695 ;
      RECT -11.165 -49.515 -11.065 -48.915 ;
      RECT -11.165 -44.575 -11.065 -44.155 ;
      RECT -11.165 -43.055 -11.065 -42.635 ;
      RECT -11.165 -38.295 -11.065 -37.695 ;
      RECT -11.165 -36.595 -11.065 -35.995 ;
      RECT -11.165 -31.655 -11.065 -31.235 ;
      RECT -11.165 -30.135 -11.065 -29.715 ;
      RECT -11.165 -25.375 -11.065 -24.775 ;
      RECT -11.165 -23.675 -11.065 -23.075 ;
      RECT -11.165 -18.735 -11.065 -18.315 ;
      RECT -11.165 -17.215 -11.065 -16.795 ;
      RECT -11.165 -12.455 -11.065 -11.855 ;
      RECT -11.165 -10.755 -11.065 -10.155 ;
      RECT -11.165 -5.815 -11.065 -5.395 ;
      RECT -11.165 -4.295 -11.065 -3.875 ;
      RECT -11.165 0.465 -11.065 1.065 ;
      RECT -11.265 -58.955 -11.165 -58.475 ;
      RECT -11.265 -57.495 -11.165 -57.075 ;
      RECT -11.685 -44.755 -11.585 -44.155 ;
      RECT -11.685 -43.055 -11.585 -42.455 ;
      RECT -11.685 -31.835 -11.585 -31.235 ;
      RECT -11.685 -30.135 -11.585 -29.535 ;
      RECT -11.685 -18.915 -11.585 -18.315 ;
      RECT -11.685 -17.215 -11.585 -16.615 ;
      RECT -11.685 -5.995 -11.585 -5.395 ;
      RECT -11.685 -4.295 -11.585 -3.695 ;
      RECT -12.505 -47.035 -11.68 -46.935 ;
      RECT -12.505 -40.275 -11.68 -40.175 ;
      RECT -12.505 -34.115 -11.68 -34.015 ;
      RECT -12.505 -27.355 -11.68 -27.255 ;
      RECT -12.505 -21.195 -11.68 -21.095 ;
      RECT -12.505 -14.435 -11.68 -14.335 ;
      RECT -12.505 -8.275 -11.68 -8.175 ;
      RECT -12.505 -1.515 -11.68 -1.415 ;
      RECT -11.865 -58.955 -11.765 -58.475 ;
      RECT -11.865 -57.495 -11.765 -57.075 ;
      RECT -11.945 -44.755 -11.845 -44.155 ;
      RECT -11.945 -43.055 -11.845 -42.455 ;
      RECT -11.945 -31.835 -11.845 -31.235 ;
      RECT -11.945 -30.135 -11.845 -29.535 ;
      RECT -11.945 -18.915 -11.845 -18.315 ;
      RECT -11.945 -17.215 -11.845 -16.615 ;
      RECT -11.945 -5.995 -11.845 -5.395 ;
      RECT -11.945 -4.295 -11.845 -3.695 ;
      RECT -12.465 -49.515 -12.365 -48.915 ;
      RECT -12.465 -44.575 -12.365 -44.155 ;
      RECT -12.465 -43.055 -12.365 -42.635 ;
      RECT -12.465 -38.295 -12.365 -37.695 ;
      RECT -12.465 -36.595 -12.365 -35.995 ;
      RECT -12.465 -31.655 -12.365 -31.235 ;
      RECT -12.465 -30.135 -12.365 -29.715 ;
      RECT -12.465 -25.375 -12.365 -24.775 ;
      RECT -12.465 -23.675 -12.365 -23.075 ;
      RECT -12.465 -18.735 -12.365 -18.315 ;
      RECT -12.465 -17.215 -12.365 -16.795 ;
      RECT -12.465 -12.455 -12.365 -11.855 ;
      RECT -12.465 -10.755 -12.365 -10.155 ;
      RECT -12.465 -5.815 -12.365 -5.395 ;
      RECT -12.465 -4.295 -12.365 -3.875 ;
      RECT -12.465 0.465 -12.365 1.065 ;
      RECT -12.985 -44.755 -12.885 -44.155 ;
      RECT -12.985 -43.055 -12.885 -42.455 ;
      RECT -12.985 -31.835 -12.885 -31.235 ;
      RECT -12.985 -30.135 -12.885 -29.535 ;
      RECT -12.985 -18.915 -12.885 -18.315 ;
      RECT -12.985 -17.215 -12.885 -16.615 ;
      RECT -12.985 -5.995 -12.885 -5.395 ;
      RECT -12.985 -4.295 -12.885 -3.695 ;
      RECT -13.805 -46.815 -12.98 -46.715 ;
      RECT -13.805 -40.495 -12.98 -40.395 ;
      RECT -13.805 -33.895 -12.98 -33.795 ;
      RECT -13.805 -27.575 -12.98 -27.475 ;
      RECT -13.805 -20.975 -12.98 -20.875 ;
      RECT -13.805 -14.655 -12.98 -14.555 ;
      RECT -13.805 -8.055 -12.98 -7.955 ;
      RECT -13.805 -1.735 -12.98 -1.635 ;
      RECT -13.245 -44.755 -13.145 -44.155 ;
      RECT -13.245 -43.055 -13.145 -42.455 ;
      RECT -13.245 -31.835 -13.145 -31.235 ;
      RECT -13.245 -30.135 -13.145 -29.535 ;
      RECT -13.245 -18.915 -13.145 -18.315 ;
      RECT -13.245 -17.215 -13.145 -16.615 ;
      RECT -13.245 -5.995 -13.145 -5.395 ;
      RECT -13.245 -4.295 -13.145 -3.695 ;
      RECT -15.105 -47.035 -13.24 -46.935 ;
      RECT -15.105 -40.275 -13.24 -40.175 ;
      RECT -15.105 -34.115 -13.24 -34.015 ;
      RECT -15.105 -27.355 -13.24 -27.255 ;
      RECT -15.105 -21.195 -13.24 -21.095 ;
      RECT -15.105 -14.435 -13.24 -14.335 ;
      RECT -15.105 -8.275 -13.24 -8.175 ;
      RECT -15.105 -1.515 -13.24 -1.415 ;
      RECT -13.765 -49.515 -13.665 -48.915 ;
      RECT -13.765 -44.575 -13.665 -44.155 ;
      RECT -13.765 -43.055 -13.665 -42.635 ;
      RECT -13.765 -38.295 -13.665 -37.695 ;
      RECT -13.765 -36.595 -13.665 -35.995 ;
      RECT -13.765 -31.655 -13.665 -31.235 ;
      RECT -13.765 -30.135 -13.665 -29.715 ;
      RECT -13.765 -25.375 -13.665 -24.775 ;
      RECT -13.765 -23.675 -13.665 -23.075 ;
      RECT -13.765 -18.735 -13.665 -18.315 ;
      RECT -13.765 -17.215 -13.665 -16.795 ;
      RECT -13.765 -12.455 -13.665 -11.855 ;
      RECT -13.765 -10.755 -13.665 -10.155 ;
      RECT -13.765 -5.815 -13.665 -5.395 ;
      RECT -13.765 -4.295 -13.665 -3.875 ;
      RECT -13.765 0.465 -13.665 1.065 ;
      RECT -14.285 -44.755 -14.185 -44.155 ;
      RECT -14.285 -43.055 -14.185 -42.455 ;
      RECT -14.285 -31.835 -14.185 -31.235 ;
      RECT -14.285 -30.135 -14.185 -29.535 ;
      RECT -14.285 -18.915 -14.185 -18.315 ;
      RECT -14.285 -17.215 -14.185 -16.615 ;
      RECT -14.285 -5.995 -14.185 -5.395 ;
      RECT -14.285 -4.295 -14.185 -3.695 ;
      RECT -14.545 -44.755 -14.445 -44.155 ;
      RECT -14.545 -43.055 -14.445 -42.455 ;
      RECT -14.545 -31.835 -14.445 -31.235 ;
      RECT -14.545 -30.135 -14.445 -29.535 ;
      RECT -14.545 -18.915 -14.445 -18.315 ;
      RECT -14.545 -17.215 -14.445 -16.615 ;
      RECT -14.545 -5.995 -14.445 -5.395 ;
      RECT -14.545 -4.295 -14.445 -3.695 ;
      RECT -15.065 -49.515 -14.965 -48.915 ;
      RECT -15.065 -44.575 -14.965 -44.155 ;
      RECT -15.065 -43.055 -14.965 -42.635 ;
      RECT -15.065 -38.295 -14.965 -37.695 ;
      RECT -15.065 -36.595 -14.965 -35.995 ;
      RECT -15.065 -31.655 -14.965 -31.235 ;
      RECT -15.065 -30.135 -14.965 -29.715 ;
      RECT -15.065 -25.375 -14.965 -24.775 ;
      RECT -15.065 -23.675 -14.965 -23.075 ;
      RECT -15.065 -18.735 -14.965 -18.315 ;
      RECT -15.065 -17.215 -14.965 -16.795 ;
      RECT -15.065 -12.455 -14.965 -11.855 ;
      RECT -15.065 -10.755 -14.965 -10.155 ;
      RECT -15.065 -5.815 -14.965 -5.395 ;
      RECT -15.065 -4.295 -14.965 -3.875 ;
      RECT -15.065 0.465 -14.965 1.065 ;
      RECT -15.585 -44.755 -15.485 -44.155 ;
      RECT -15.585 -43.055 -15.485 -42.455 ;
      RECT -15.585 -31.835 -15.485 -31.235 ;
      RECT -15.585 -30.135 -15.485 -29.535 ;
      RECT -15.585 -18.915 -15.485 -18.315 ;
      RECT -15.585 -17.215 -15.485 -16.615 ;
      RECT -15.585 -5.995 -15.485 -5.395 ;
      RECT -15.585 -4.295 -15.485 -3.695 ;
      RECT -15.845 -44.755 -15.745 -44.155 ;
      RECT -15.845 -43.055 -15.745 -42.455 ;
      RECT -15.845 -31.835 -15.745 -31.235 ;
      RECT -15.845 -30.135 -15.745 -29.535 ;
      RECT -15.845 -18.915 -15.745 -18.315 ;
      RECT -15.845 -17.215 -15.745 -16.615 ;
      RECT -15.845 -5.995 -15.745 -5.395 ;
      RECT -15.845 -4.295 -15.745 -3.695 ;
      RECT -29.865 -48.575 -15.84 -48.475 ;
      RECT -29.865 -38.735 -15.84 -38.635 ;
      RECT -29.865 -35.655 -15.84 -35.555 ;
      RECT -29.865 -25.815 -15.84 -25.715 ;
      RECT -29.865 -22.735 -15.84 -22.635 ;
      RECT -29.865 -12.895 -15.84 -12.795 ;
      RECT -29.865 -9.815 -15.84 -9.715 ;
      RECT -29.865 0.025 -15.84 0.125 ;
      RECT -16.365 -49.515 -16.265 -48.915 ;
      RECT -16.365 -44.575 -16.265 -44.155 ;
      RECT -16.365 -43.055 -16.265 -42.635 ;
      RECT -16.365 -38.295 -16.265 -37.695 ;
      RECT -16.365 -36.595 -16.265 -35.995 ;
      RECT -16.365 -31.655 -16.265 -31.235 ;
      RECT -16.365 -30.135 -16.265 -29.715 ;
      RECT -16.365 -25.375 -16.265 -24.775 ;
      RECT -16.365 -23.675 -16.265 -23.075 ;
      RECT -16.365 -18.735 -16.265 -18.315 ;
      RECT -16.365 -17.215 -16.265 -16.795 ;
      RECT -16.365 -12.455 -16.265 -11.855 ;
      RECT -16.365 -10.755 -16.265 -10.155 ;
      RECT -16.365 -5.815 -16.265 -5.395 ;
      RECT -16.365 -4.295 -16.265 -3.875 ;
      RECT -16.365 0.465 -16.265 1.065 ;
      RECT -16.885 -44.755 -16.785 -44.155 ;
      RECT -16.885 -43.055 -16.785 -42.455 ;
      RECT -16.885 -31.835 -16.785 -31.235 ;
      RECT -16.885 -30.135 -16.785 -29.535 ;
      RECT -16.885 -18.915 -16.785 -18.315 ;
      RECT -16.885 -17.215 -16.785 -16.615 ;
      RECT -16.885 -5.995 -16.785 -5.395 ;
      RECT -16.885 -4.295 -16.785 -3.695 ;
      RECT -17.705 -47.035 -16.88 -46.935 ;
      RECT -17.705 -40.275 -16.88 -40.175 ;
      RECT -17.705 -34.115 -16.88 -34.015 ;
      RECT -17.705 -27.355 -16.88 -27.255 ;
      RECT -17.705 -21.195 -16.88 -21.095 ;
      RECT -17.705 -14.435 -16.88 -14.335 ;
      RECT -17.705 -8.275 -16.88 -8.175 ;
      RECT -17.705 -1.515 -16.88 -1.415 ;
      RECT -17.145 -44.755 -17.045 -44.155 ;
      RECT -17.145 -43.055 -17.045 -42.455 ;
      RECT -17.145 -31.835 -17.045 -31.235 ;
      RECT -17.145 -30.135 -17.045 -29.535 ;
      RECT -17.145 -18.915 -17.045 -18.315 ;
      RECT -17.145 -17.215 -17.045 -16.615 ;
      RECT -17.145 -5.995 -17.045 -5.395 ;
      RECT -17.145 -4.295 -17.045 -3.695 ;
      RECT -17.665 -49.515 -17.565 -48.915 ;
      RECT -17.665 -44.575 -17.565 -44.155 ;
      RECT -17.665 -43.055 -17.565 -42.635 ;
      RECT -17.665 -38.295 -17.565 -37.695 ;
      RECT -17.665 -36.595 -17.565 -35.995 ;
      RECT -17.665 -31.655 -17.565 -31.235 ;
      RECT -17.665 -30.135 -17.565 -29.715 ;
      RECT -17.665 -25.375 -17.565 -24.775 ;
      RECT -17.665 -23.675 -17.565 -23.075 ;
      RECT -17.665 -18.735 -17.565 -18.315 ;
      RECT -17.665 -17.215 -17.565 -16.795 ;
      RECT -17.665 -12.455 -17.565 -11.855 ;
      RECT -17.665 -10.755 -17.565 -10.155 ;
      RECT -17.665 -5.815 -17.565 -5.395 ;
      RECT -17.665 -4.295 -17.565 -3.875 ;
      RECT -17.665 0.465 -17.565 1.065 ;
      RECT -18.185 -44.755 -18.085 -44.155 ;
      RECT -18.185 -43.055 -18.085 -42.455 ;
      RECT -18.185 -31.835 -18.085 -31.235 ;
      RECT -18.185 -30.135 -18.085 -29.535 ;
      RECT -18.185 -18.915 -18.085 -18.315 ;
      RECT -18.185 -17.215 -18.085 -16.615 ;
      RECT -18.185 -5.995 -18.085 -5.395 ;
      RECT -18.185 -4.295 -18.085 -3.695 ;
      RECT -19.005 -46.815 -18.18 -46.715 ;
      RECT -19.005 -40.495 -18.18 -40.395 ;
      RECT -19.005 -33.895 -18.18 -33.795 ;
      RECT -19.005 -27.575 -18.18 -27.475 ;
      RECT -19.005 -20.975 -18.18 -20.875 ;
      RECT -19.005 -14.655 -18.18 -14.555 ;
      RECT -19.005 -8.055 -18.18 -7.955 ;
      RECT -19.005 -1.735 -18.18 -1.635 ;
      RECT -18.445 -44.755 -18.345 -44.155 ;
      RECT -18.445 -43.055 -18.345 -42.455 ;
      RECT -18.445 -31.835 -18.345 -31.235 ;
      RECT -18.445 -30.135 -18.345 -29.535 ;
      RECT -18.445 -18.915 -18.345 -18.315 ;
      RECT -18.445 -17.215 -18.345 -16.615 ;
      RECT -18.445 -5.995 -18.345 -5.395 ;
      RECT -18.445 -4.295 -18.345 -3.695 ;
      RECT -20.305 -47.035 -18.44 -46.935 ;
      RECT -20.305 -40.275 -18.44 -40.175 ;
      RECT -20.305 -34.115 -18.44 -34.015 ;
      RECT -20.305 -27.355 -18.44 -27.255 ;
      RECT -20.305 -21.195 -18.44 -21.095 ;
      RECT -20.305 -14.435 -18.44 -14.335 ;
      RECT -20.305 -8.275 -18.44 -8.175 ;
      RECT -20.305 -1.515 -18.44 -1.415 ;
      RECT -18.965 -49.515 -18.865 -48.915 ;
      RECT -18.965 -44.575 -18.865 -44.155 ;
      RECT -18.965 -43.055 -18.865 -42.635 ;
      RECT -18.965 -38.295 -18.865 -37.695 ;
      RECT -18.965 -36.595 -18.865 -35.995 ;
      RECT -18.965 -31.655 -18.865 -31.235 ;
      RECT -18.965 -30.135 -18.865 -29.715 ;
      RECT -18.965 -25.375 -18.865 -24.775 ;
      RECT -18.965 -23.675 -18.865 -23.075 ;
      RECT -18.965 -18.735 -18.865 -18.315 ;
      RECT -18.965 -17.215 -18.865 -16.795 ;
      RECT -18.965 -12.455 -18.865 -11.855 ;
      RECT -18.965 -10.755 -18.865 -10.155 ;
      RECT -18.965 -5.815 -18.865 -5.395 ;
      RECT -18.965 -4.295 -18.865 -3.875 ;
      RECT -18.965 0.465 -18.865 1.065 ;
      RECT -19.485 -44.755 -19.385 -44.155 ;
      RECT -19.485 -43.055 -19.385 -42.455 ;
      RECT -19.485 -31.835 -19.385 -31.235 ;
      RECT -19.485 -30.135 -19.385 -29.535 ;
      RECT -19.485 -18.915 -19.385 -18.315 ;
      RECT -19.485 -17.215 -19.385 -16.615 ;
      RECT -19.485 -5.995 -19.385 -5.395 ;
      RECT -19.485 -4.295 -19.385 -3.695 ;
      RECT -19.745 -44.755 -19.645 -44.155 ;
      RECT -19.745 -43.055 -19.645 -42.455 ;
      RECT -19.745 -31.835 -19.645 -31.235 ;
      RECT -19.745 -30.135 -19.645 -29.535 ;
      RECT -19.745 -18.915 -19.645 -18.315 ;
      RECT -19.745 -17.215 -19.645 -16.615 ;
      RECT -19.745 -5.995 -19.645 -5.395 ;
      RECT -19.745 -4.295 -19.645 -3.695 ;
      RECT -20.265 -49.515 -20.165 -48.915 ;
      RECT -20.265 -44.575 -20.165 -44.155 ;
      RECT -20.265 -43.055 -20.165 -42.635 ;
      RECT -20.265 -38.295 -20.165 -37.695 ;
      RECT -20.265 -36.595 -20.165 -35.995 ;
      RECT -20.265 -31.655 -20.165 -31.235 ;
      RECT -20.265 -30.135 -20.165 -29.715 ;
      RECT -20.265 -25.375 -20.165 -24.775 ;
      RECT -20.265 -23.675 -20.165 -23.075 ;
      RECT -20.265 -18.735 -20.165 -18.315 ;
      RECT -20.265 -17.215 -20.165 -16.795 ;
      RECT -20.265 -12.455 -20.165 -11.855 ;
      RECT -20.265 -10.755 -20.165 -10.155 ;
      RECT -20.265 -5.815 -20.165 -5.395 ;
      RECT -20.265 -4.295 -20.165 -3.875 ;
      RECT -20.265 0.465 -20.165 1.065 ;
      RECT -20.785 -44.755 -20.685 -44.155 ;
      RECT -20.785 -43.055 -20.685 -42.455 ;
      RECT -20.785 -31.835 -20.685 -31.235 ;
      RECT -20.785 -30.135 -20.685 -29.535 ;
      RECT -20.785 -18.915 -20.685 -18.315 ;
      RECT -20.785 -17.215 -20.685 -16.615 ;
      RECT -20.785 -5.995 -20.685 -5.395 ;
      RECT -20.785 -4.295 -20.685 -3.695 ;
      RECT -29.865 -48.135 -20.78 -48.035 ;
      RECT -29.865 -39.175 -20.78 -39.075 ;
      RECT -29.865 -35.215 -20.78 -35.115 ;
      RECT -29.865 -26.255 -20.78 -26.155 ;
      RECT -29.865 -22.295 -20.78 -22.195 ;
      RECT -29.865 -13.335 -20.78 -13.235 ;
      RECT -29.865 -9.375 -20.78 -9.275 ;
      RECT -29.865 -0.415 -20.78 -0.315 ;
      RECT -21.045 -44.755 -20.945 -44.155 ;
      RECT -21.045 -43.055 -20.945 -42.455 ;
      RECT -21.045 -31.835 -20.945 -31.235 ;
      RECT -21.045 -30.135 -20.945 -29.535 ;
      RECT -21.045 -18.915 -20.945 -18.315 ;
      RECT -21.045 -17.215 -20.945 -16.615 ;
      RECT -21.045 -5.995 -20.945 -5.395 ;
      RECT -21.045 -4.295 -20.945 -3.695 ;
      RECT -21.565 -49.515 -21.465 -48.915 ;
      RECT -21.565 -44.575 -21.465 -44.155 ;
      RECT -21.565 -43.055 -21.465 -42.635 ;
      RECT -21.565 -38.295 -21.465 -37.695 ;
      RECT -21.565 -36.595 -21.465 -35.995 ;
      RECT -21.565 -31.655 -21.465 -31.235 ;
      RECT -21.565 -30.135 -21.465 -29.715 ;
      RECT -21.565 -25.375 -21.465 -24.775 ;
      RECT -21.565 -23.675 -21.465 -23.075 ;
      RECT -21.565 -18.735 -21.465 -18.315 ;
      RECT -21.565 -17.215 -21.465 -16.795 ;
      RECT -21.565 -12.455 -21.465 -11.855 ;
      RECT -21.565 -10.755 -21.465 -10.155 ;
      RECT -21.565 -5.815 -21.465 -5.395 ;
      RECT -21.565 -4.295 -21.465 -3.875 ;
      RECT -21.565 0.465 -21.465 1.065 ;
      RECT -22.085 -44.755 -21.985 -44.155 ;
      RECT -22.085 -43.055 -21.985 -42.455 ;
      RECT -22.085 -31.835 -21.985 -31.235 ;
      RECT -22.085 -30.135 -21.985 -29.535 ;
      RECT -22.085 -18.915 -21.985 -18.315 ;
      RECT -22.085 -17.215 -21.985 -16.615 ;
      RECT -22.085 -5.995 -21.985 -5.395 ;
      RECT -22.085 -4.295 -21.985 -3.695 ;
      RECT -22.905 -47.035 -22.08 -46.935 ;
      RECT -22.905 -40.275 -22.08 -40.175 ;
      RECT -22.905 -34.115 -22.08 -34.015 ;
      RECT -22.905 -27.355 -22.08 -27.255 ;
      RECT -22.905 -21.195 -22.08 -21.095 ;
      RECT -22.905 -14.435 -22.08 -14.335 ;
      RECT -22.905 -8.275 -22.08 -8.175 ;
      RECT -22.905 -1.515 -22.08 -1.415 ;
      RECT -22.345 -44.755 -22.245 -44.155 ;
      RECT -22.345 -43.055 -22.245 -42.455 ;
      RECT -22.345 -31.835 -22.245 -31.235 ;
      RECT -22.345 -30.135 -22.245 -29.535 ;
      RECT -22.345 -18.915 -22.245 -18.315 ;
      RECT -22.345 -17.215 -22.245 -16.615 ;
      RECT -22.345 -5.995 -22.245 -5.395 ;
      RECT -22.345 -4.295 -22.245 -3.695 ;
      RECT -22.865 -49.515 -22.765 -48.915 ;
      RECT -22.865 -44.575 -22.765 -44.155 ;
      RECT -22.865 -43.055 -22.765 -42.635 ;
      RECT -22.865 -38.295 -22.765 -37.695 ;
      RECT -22.865 -36.595 -22.765 -35.995 ;
      RECT -22.865 -31.655 -22.765 -31.235 ;
      RECT -22.865 -30.135 -22.765 -29.715 ;
      RECT -22.865 -25.375 -22.765 -24.775 ;
      RECT -22.865 -23.675 -22.765 -23.075 ;
      RECT -22.865 -18.735 -22.765 -18.315 ;
      RECT -22.865 -17.215 -22.765 -16.795 ;
      RECT -22.865 -12.455 -22.765 -11.855 ;
      RECT -22.865 -10.755 -22.765 -10.155 ;
      RECT -22.865 -5.815 -22.765 -5.395 ;
      RECT -22.865 -4.295 -22.765 -3.875 ;
      RECT -22.865 0.465 -22.765 1.065 ;
      RECT -23.385 -44.755 -23.285 -44.155 ;
      RECT -23.385 -43.055 -23.285 -42.455 ;
      RECT -23.385 -31.835 -23.285 -31.235 ;
      RECT -23.385 -30.135 -23.285 -29.535 ;
      RECT -23.385 -18.915 -23.285 -18.315 ;
      RECT -23.385 -17.215 -23.285 -16.615 ;
      RECT -23.385 -5.995 -23.285 -5.395 ;
      RECT -23.385 -4.295 -23.285 -3.695 ;
      RECT -24.205 -46.815 -23.38 -46.715 ;
      RECT -24.205 -40.495 -23.38 -40.395 ;
      RECT -24.205 -33.895 -23.38 -33.795 ;
      RECT -24.205 -27.575 -23.38 -27.475 ;
      RECT -24.205 -20.975 -23.38 -20.875 ;
      RECT -24.205 -14.655 -23.38 -14.555 ;
      RECT -24.205 -8.055 -23.38 -7.955 ;
      RECT -24.205 -1.735 -23.38 -1.635 ;
      RECT -23.645 -44.755 -23.545 -44.155 ;
      RECT -23.645 -43.055 -23.545 -42.455 ;
      RECT -23.645 -31.835 -23.545 -31.235 ;
      RECT -23.645 -30.135 -23.545 -29.535 ;
      RECT -23.645 -18.915 -23.545 -18.315 ;
      RECT -23.645 -17.215 -23.545 -16.615 ;
      RECT -23.645 -5.995 -23.545 -5.395 ;
      RECT -23.645 -4.295 -23.545 -3.695 ;
      RECT -25.505 -47.035 -23.64 -46.935 ;
      RECT -25.505 -40.275 -23.64 -40.175 ;
      RECT -25.505 -34.115 -23.64 -34.015 ;
      RECT -25.505 -27.355 -23.64 -27.255 ;
      RECT -25.505 -21.195 -23.64 -21.095 ;
      RECT -25.505 -14.435 -23.64 -14.335 ;
      RECT -25.505 -8.275 -23.64 -8.175 ;
      RECT -25.505 -1.515 -23.64 -1.415 ;
      RECT -24.165 -49.515 -24.065 -48.915 ;
      RECT -24.165 -44.575 -24.065 -44.155 ;
      RECT -24.165 -43.055 -24.065 -42.635 ;
      RECT -24.165 -38.295 -24.065 -37.695 ;
      RECT -24.165 -36.595 -24.065 -35.995 ;
      RECT -24.165 -31.655 -24.065 -31.235 ;
      RECT -24.165 -30.135 -24.065 -29.715 ;
      RECT -24.165 -25.375 -24.065 -24.775 ;
      RECT -24.165 -23.675 -24.065 -23.075 ;
      RECT -24.165 -18.735 -24.065 -18.315 ;
      RECT -24.165 -17.215 -24.065 -16.795 ;
      RECT -24.165 -12.455 -24.065 -11.855 ;
      RECT -24.165 -10.755 -24.065 -10.155 ;
      RECT -24.165 -5.815 -24.065 -5.395 ;
      RECT -24.165 -4.295 -24.065 -3.875 ;
      RECT -24.165 0.465 -24.065 1.065 ;
      RECT -24.685 -44.755 -24.585 -44.155 ;
      RECT -24.685 -43.055 -24.585 -42.455 ;
      RECT -24.685 -31.835 -24.585 -31.235 ;
      RECT -24.685 -30.135 -24.585 -29.535 ;
      RECT -24.685 -18.915 -24.585 -18.315 ;
      RECT -24.685 -17.215 -24.585 -16.615 ;
      RECT -24.685 -5.995 -24.585 -5.395 ;
      RECT -24.685 -4.295 -24.585 -3.695 ;
      RECT -24.945 -44.755 -24.845 -44.155 ;
      RECT -24.945 -43.055 -24.845 -42.455 ;
      RECT -24.945 -31.835 -24.845 -31.235 ;
      RECT -24.945 -30.135 -24.845 -29.535 ;
      RECT -24.945 -18.915 -24.845 -18.315 ;
      RECT -24.945 -17.215 -24.845 -16.615 ;
      RECT -24.945 -5.995 -24.845 -5.395 ;
      RECT -24.945 -4.295 -24.845 -3.695 ;
      RECT -25.465 -49.515 -25.365 -48.915 ;
      RECT -25.465 -44.575 -25.365 -44.155 ;
      RECT -25.465 -43.055 -25.365 -42.635 ;
      RECT -25.465 -38.295 -25.365 -37.695 ;
      RECT -25.465 -36.595 -25.365 -35.995 ;
      RECT -25.465 -31.655 -25.365 -31.235 ;
      RECT -25.465 -30.135 -25.365 -29.715 ;
      RECT -25.465 -25.375 -25.365 -24.775 ;
      RECT -25.465 -23.675 -25.365 -23.075 ;
      RECT -25.465 -18.735 -25.365 -18.315 ;
      RECT -25.465 -17.215 -25.365 -16.795 ;
      RECT -25.465 -12.455 -25.365 -11.855 ;
      RECT -25.465 -10.755 -25.365 -10.155 ;
      RECT -25.465 -5.815 -25.365 -5.395 ;
      RECT -25.465 -4.295 -25.365 -3.875 ;
      RECT -25.465 0.465 -25.365 1.065 ;
      RECT -25.985 -44.755 -25.885 -44.155 ;
      RECT -25.985 -43.055 -25.885 -42.455 ;
      RECT -25.985 -31.835 -25.885 -31.235 ;
      RECT -25.985 -30.135 -25.885 -29.535 ;
      RECT -25.985 -18.915 -25.885 -18.315 ;
      RECT -25.985 -17.215 -25.885 -16.615 ;
      RECT -25.985 -5.995 -25.885 -5.395 ;
      RECT -25.985 -4.295 -25.885 -3.695 ;
      RECT -26.245 -44.755 -26.145 -44.155 ;
      RECT -26.245 -43.055 -26.145 -42.455 ;
      RECT -26.245 -31.835 -26.145 -31.235 ;
      RECT -26.245 -30.135 -26.145 -29.535 ;
      RECT -26.245 -18.915 -26.145 -18.315 ;
      RECT -26.245 -17.215 -26.145 -16.615 ;
      RECT -26.245 -5.995 -26.145 -5.395 ;
      RECT -26.245 -4.295 -26.145 -3.695 ;
      RECT -26.865 2.165 -26.765 2.645 ;
      RECT -26.865 4.645 -26.765 5.065 ;
      RECT -27.465 2.165 -27.365 2.645 ;
      RECT -27.465 4.645 -27.365 5.065 ;
      RECT -28.065 2.165 -27.965 2.645 ;
      RECT -28.065 4.645 -27.965 5.065 ;
      RECT -28.665 2.165 -28.565 2.645 ;
      RECT -28.665 4.645 -28.565 5.065 ;
      RECT -29.265 2.165 -29.165 2.645 ;
      RECT -29.265 4.645 -29.165 5.065 ;
    LAYER V1 ;
      RECT 38.275 -57.245 38.375 -57.145 ;
      RECT 38.275 -53.195 38.375 -53.095 ;
      RECT 38.275 -52.955 38.375 -52.855 ;
      RECT 38.275 -52.715 38.375 -52.615 ;
      RECT 38.275 -52.475 38.375 -52.375 ;
      RECT 38.015 -53.195 38.115 -53.095 ;
      RECT 38.015 -52.955 38.115 -52.855 ;
      RECT 38.015 -52.715 38.115 -52.615 ;
      RECT 38.015 -52.475 38.115 -52.375 ;
      RECT 38.015 -48.5 38.115 -48.4 ;
      RECT 38.015 -45.27 38.115 -45.17 ;
      RECT 38.015 -42.04 38.115 -41.94 ;
      RECT 38.015 -38.81 38.115 -38.71 ;
      RECT 38.015 -35.58 38.115 -35.48 ;
      RECT 38.015 -32.35 38.115 -32.25 ;
      RECT 38.015 -29.12 38.115 -29.02 ;
      RECT 38.015 -25.89 38.115 -25.79 ;
      RECT 38.015 -22.66 38.115 -22.56 ;
      RECT 38.015 -19.43 38.115 -19.33 ;
      RECT 38.015 -16.2 38.115 -16.1 ;
      RECT 38.015 -12.97 38.115 -12.87 ;
      RECT 38.015 -9.74 38.115 -9.64 ;
      RECT 38.015 -6.51 38.115 -6.41 ;
      RECT 38.015 -3.28 38.115 -3.18 ;
      RECT 38.015 -0.05 38.115 0.05 ;
      RECT 38.015 2.245 38.115 2.345 ;
      RECT 38.015 2.485 38.115 2.585 ;
      RECT 38.015 2.725 38.115 2.825 ;
      RECT 38.015 2.965 38.115 3.065 ;
      RECT 37.725 -60.485 37.825 -60.385 ;
      RECT 37.725 -60.285 37.825 -60.185 ;
      RECT 37.725 -59.015 37.825 -58.915 ;
      RECT 37.585 -53.195 37.685 -53.095 ;
      RECT 37.585 -52.955 37.685 -52.855 ;
      RECT 37.585 -52.715 37.685 -52.615 ;
      RECT 37.585 -52.475 37.685 -52.375 ;
      RECT 37.585 -48.5 37.685 -48.4 ;
      RECT 37.585 -45.27 37.685 -45.17 ;
      RECT 37.585 -42.04 37.685 -41.94 ;
      RECT 37.585 -38.81 37.685 -38.71 ;
      RECT 37.585 -35.58 37.685 -35.48 ;
      RECT 37.585 -32.35 37.685 -32.25 ;
      RECT 37.585 -29.12 37.685 -29.02 ;
      RECT 37.585 -25.89 37.685 -25.79 ;
      RECT 37.585 -22.66 37.685 -22.56 ;
      RECT 37.585 -19.43 37.685 -19.33 ;
      RECT 37.585 -16.2 37.685 -16.1 ;
      RECT 37.585 -12.97 37.685 -12.87 ;
      RECT 37.585 -9.74 37.685 -9.64 ;
      RECT 37.585 -6.51 37.685 -6.41 ;
      RECT 37.585 -3.28 37.685 -3.18 ;
      RECT 37.585 -0.05 37.685 0.05 ;
      RECT 37.585 2.245 37.685 2.345 ;
      RECT 37.585 2.485 37.685 2.585 ;
      RECT 37.585 2.725 37.685 2.825 ;
      RECT 37.585 2.965 37.685 3.065 ;
      RECT 37.325 -56.965 37.425 -56.865 ;
      RECT 37.325 -53.195 37.425 -53.095 ;
      RECT 37.325 -52.955 37.425 -52.855 ;
      RECT 37.325 -52.715 37.425 -52.615 ;
      RECT 37.325 -52.475 37.425 -52.375 ;
      RECT 37.135 -60.265 37.235 -60.165 ;
      RECT 37.135 -60.005 37.235 -59.905 ;
      RECT 37.135 -59.03 37.235 -58.93 ;
      RECT 37.135 -58.83 37.235 -58.73 ;
      RECT 37.075 -57.245 37.175 -57.145 ;
      RECT 37.075 -53.195 37.175 -53.095 ;
      RECT 37.075 -52.955 37.175 -52.855 ;
      RECT 37.075 -52.715 37.175 -52.615 ;
      RECT 37.075 -52.475 37.175 -52.375 ;
      RECT 36.835 -57.47 36.935 -57.37 ;
      RECT 36.835 -56.965 36.935 -56.865 ;
      RECT 36.815 -53.195 36.915 -53.095 ;
      RECT 36.815 -52.955 36.915 -52.855 ;
      RECT 36.815 -52.715 36.915 -52.615 ;
      RECT 36.815 -52.475 36.915 -52.375 ;
      RECT 36.815 -48.5 36.915 -48.4 ;
      RECT 36.815 -45.27 36.915 -45.17 ;
      RECT 36.815 -42.04 36.915 -41.94 ;
      RECT 36.815 -38.81 36.915 -38.71 ;
      RECT 36.815 -35.58 36.915 -35.48 ;
      RECT 36.815 -32.35 36.915 -32.25 ;
      RECT 36.815 -29.12 36.915 -29.02 ;
      RECT 36.815 -25.89 36.915 -25.79 ;
      RECT 36.815 -22.66 36.915 -22.56 ;
      RECT 36.815 -19.43 36.915 -19.33 ;
      RECT 36.815 -16.2 36.915 -16.1 ;
      RECT 36.815 -12.97 36.915 -12.87 ;
      RECT 36.815 -9.74 36.915 -9.64 ;
      RECT 36.815 -6.51 36.915 -6.41 ;
      RECT 36.815 -3.28 36.915 -3.18 ;
      RECT 36.815 -0.05 36.915 0.05 ;
      RECT 36.815 2.245 36.915 2.345 ;
      RECT 36.815 2.485 36.915 2.585 ;
      RECT 36.815 2.725 36.915 2.825 ;
      RECT 36.815 2.965 36.915 3.065 ;
      RECT 36.565 -57.875 36.665 -57.775 ;
      RECT 36.385 -53.195 36.485 -53.095 ;
      RECT 36.385 -52.955 36.485 -52.855 ;
      RECT 36.385 -52.715 36.485 -52.615 ;
      RECT 36.385 -52.475 36.485 -52.375 ;
      RECT 36.385 -48.5 36.485 -48.4 ;
      RECT 36.385 -45.27 36.485 -45.17 ;
      RECT 36.385 -42.04 36.485 -41.94 ;
      RECT 36.385 -38.81 36.485 -38.71 ;
      RECT 36.385 -35.58 36.485 -35.48 ;
      RECT 36.385 -32.35 36.485 -32.25 ;
      RECT 36.385 -29.12 36.485 -29.02 ;
      RECT 36.385 -25.89 36.485 -25.79 ;
      RECT 36.385 -22.66 36.485 -22.56 ;
      RECT 36.385 -19.43 36.485 -19.33 ;
      RECT 36.385 -16.2 36.485 -16.1 ;
      RECT 36.385 -12.97 36.485 -12.87 ;
      RECT 36.385 -9.74 36.485 -9.64 ;
      RECT 36.385 -6.51 36.485 -6.41 ;
      RECT 36.385 -3.28 36.485 -3.18 ;
      RECT 36.385 -0.05 36.485 0.05 ;
      RECT 36.385 2.245 36.485 2.345 ;
      RECT 36.385 2.485 36.485 2.585 ;
      RECT 36.385 2.725 36.485 2.825 ;
      RECT 36.385 2.965 36.485 3.065 ;
      RECT 36.24 -57.875 36.34 -57.775 ;
      RECT 36.125 -56.965 36.225 -56.865 ;
      RECT 36.125 -53.195 36.225 -53.095 ;
      RECT 36.125 -52.955 36.225 -52.855 ;
      RECT 36.125 -52.715 36.225 -52.615 ;
      RECT 36.125 -52.475 36.225 -52.375 ;
      RECT 35.875 -57.245 35.975 -57.145 ;
      RECT 35.875 -56.425 35.975 -56.325 ;
      RECT 35.875 -56.185 35.975 -56.085 ;
      RECT 35.875 -55.945 35.975 -55.845 ;
      RECT 35.875 -55.705 35.975 -55.605 ;
      RECT 35.705 -60.485 35.805 -60.385 ;
      RECT 35.705 -60.285 35.805 -60.185 ;
      RECT 35.705 -59.015 35.805 -58.915 ;
      RECT 35.615 -56.425 35.715 -56.325 ;
      RECT 35.615 -56.185 35.715 -56.085 ;
      RECT 35.615 -55.945 35.715 -55.845 ;
      RECT 35.615 -55.705 35.715 -55.605 ;
      RECT 35.615 -48.5 35.715 -48.4 ;
      RECT 35.615 -45.27 35.715 -45.17 ;
      RECT 35.615 -42.04 35.715 -41.94 ;
      RECT 35.615 -38.81 35.715 -38.71 ;
      RECT 35.615 -35.58 35.715 -35.48 ;
      RECT 35.615 -32.35 35.715 -32.25 ;
      RECT 35.615 -29.12 35.715 -29.02 ;
      RECT 35.615 -25.89 35.715 -25.79 ;
      RECT 35.615 -22.66 35.715 -22.56 ;
      RECT 35.615 -19.43 35.715 -19.33 ;
      RECT 35.615 -16.2 35.715 -16.1 ;
      RECT 35.615 -12.97 35.715 -12.87 ;
      RECT 35.615 -9.74 35.715 -9.64 ;
      RECT 35.615 -6.51 35.715 -6.41 ;
      RECT 35.615 -3.28 35.715 -3.18 ;
      RECT 35.615 -0.05 35.715 0.05 ;
      RECT 35.615 2.245 35.715 2.345 ;
      RECT 35.615 2.485 35.715 2.585 ;
      RECT 35.615 2.725 35.715 2.825 ;
      RECT 35.615 2.965 35.715 3.065 ;
      RECT 35.185 -56.425 35.285 -56.325 ;
      RECT 35.185 -56.185 35.285 -56.085 ;
      RECT 35.185 -55.945 35.285 -55.845 ;
      RECT 35.185 -55.705 35.285 -55.605 ;
      RECT 35.185 -48.5 35.285 -48.4 ;
      RECT 35.185 -45.27 35.285 -45.17 ;
      RECT 35.185 -42.04 35.285 -41.94 ;
      RECT 35.185 -38.81 35.285 -38.71 ;
      RECT 35.185 -35.58 35.285 -35.48 ;
      RECT 35.185 -32.35 35.285 -32.25 ;
      RECT 35.185 -29.12 35.285 -29.02 ;
      RECT 35.185 -25.89 35.285 -25.79 ;
      RECT 35.185 -22.66 35.285 -22.56 ;
      RECT 35.185 -19.43 35.285 -19.33 ;
      RECT 35.185 -16.2 35.285 -16.1 ;
      RECT 35.185 -12.97 35.285 -12.87 ;
      RECT 35.185 -9.74 35.285 -9.64 ;
      RECT 35.185 -6.51 35.285 -6.41 ;
      RECT 35.185 -3.28 35.285 -3.18 ;
      RECT 35.185 -0.05 35.285 0.05 ;
      RECT 35.185 2.245 35.285 2.345 ;
      RECT 35.185 2.485 35.285 2.585 ;
      RECT 35.185 2.725 35.285 2.825 ;
      RECT 35.185 2.965 35.285 3.065 ;
      RECT 35.115 -60.265 35.215 -60.165 ;
      RECT 35.115 -60.005 35.215 -59.905 ;
      RECT 35.115 -59.045 35.215 -58.945 ;
      RECT 35.115 -58.845 35.215 -58.745 ;
      RECT 34.925 -56.965 35.025 -56.865 ;
      RECT 34.925 -56.425 35.025 -56.325 ;
      RECT 34.925 -56.185 35.025 -56.085 ;
      RECT 34.925 -55.945 35.025 -55.845 ;
      RECT 34.925 -55.705 35.025 -55.605 ;
      RECT 34.675 -57.245 34.775 -57.145 ;
      RECT 34.675 -56.425 34.775 -56.325 ;
      RECT 34.675 -56.185 34.775 -56.085 ;
      RECT 34.675 -55.945 34.775 -55.845 ;
      RECT 34.675 -55.705 34.775 -55.605 ;
      RECT 34.415 -56.425 34.515 -56.325 ;
      RECT 34.415 -56.185 34.515 -56.085 ;
      RECT 34.415 -55.945 34.515 -55.845 ;
      RECT 34.415 -55.705 34.515 -55.605 ;
      RECT 34.415 -48.5 34.515 -48.4 ;
      RECT 34.415 -45.27 34.515 -45.17 ;
      RECT 34.415 -42.04 34.515 -41.94 ;
      RECT 34.415 -38.81 34.515 -38.71 ;
      RECT 34.415 -35.58 34.515 -35.48 ;
      RECT 34.415 -32.35 34.515 -32.25 ;
      RECT 34.415 -29.12 34.515 -29.02 ;
      RECT 34.415 -25.89 34.515 -25.79 ;
      RECT 34.415 -22.66 34.515 -22.56 ;
      RECT 34.415 -19.43 34.515 -19.33 ;
      RECT 34.415 -16.2 34.515 -16.1 ;
      RECT 34.415 -12.97 34.515 -12.87 ;
      RECT 34.415 -9.74 34.515 -9.64 ;
      RECT 34.415 -6.51 34.515 -6.41 ;
      RECT 34.415 -3.28 34.515 -3.18 ;
      RECT 34.415 -0.05 34.515 0.05 ;
      RECT 34.415 2.245 34.515 2.345 ;
      RECT 34.415 2.485 34.515 2.585 ;
      RECT 34.415 2.725 34.515 2.825 ;
      RECT 34.415 2.965 34.515 3.065 ;
      RECT 34.315 -61.745 34.415 -61.645 ;
      RECT 34.315 -61.545 34.415 -61.445 ;
      RECT 33.985 -56.425 34.085 -56.325 ;
      RECT 33.985 -56.185 34.085 -56.085 ;
      RECT 33.985 -55.945 34.085 -55.845 ;
      RECT 33.985 -55.705 34.085 -55.605 ;
      RECT 33.985 -48.5 34.085 -48.4 ;
      RECT 33.985 -45.27 34.085 -45.17 ;
      RECT 33.985 -42.04 34.085 -41.94 ;
      RECT 33.985 -38.81 34.085 -38.71 ;
      RECT 33.985 -35.58 34.085 -35.48 ;
      RECT 33.985 -32.35 34.085 -32.25 ;
      RECT 33.985 -29.12 34.085 -29.02 ;
      RECT 33.985 -25.89 34.085 -25.79 ;
      RECT 33.985 -22.66 34.085 -22.56 ;
      RECT 33.985 -19.43 34.085 -19.33 ;
      RECT 33.985 -16.2 34.085 -16.1 ;
      RECT 33.985 -12.97 34.085 -12.87 ;
      RECT 33.985 -9.74 34.085 -9.64 ;
      RECT 33.985 -6.51 34.085 -6.41 ;
      RECT 33.985 -3.28 34.085 -3.18 ;
      RECT 33.985 -0.05 34.085 0.05 ;
      RECT 33.985 2.245 34.085 2.345 ;
      RECT 33.985 2.485 34.085 2.585 ;
      RECT 33.985 2.725 34.085 2.825 ;
      RECT 33.985 2.965 34.085 3.065 ;
      RECT 33.965 -60.265 34.065 -60.165 ;
      RECT 33.965 -59.815 34.065 -59.715 ;
      RECT 33.965 -59.015 34.065 -58.915 ;
      RECT 33.725 -61.745 33.825 -61.645 ;
      RECT 33.725 -61.545 33.825 -61.445 ;
      RECT 33.725 -56.965 33.825 -56.865 ;
      RECT 33.725 -56.425 33.825 -56.325 ;
      RECT 33.725 -56.185 33.825 -56.085 ;
      RECT 33.725 -55.945 33.825 -55.845 ;
      RECT 33.725 -55.705 33.825 -55.605 ;
      RECT 33.475 -57.245 33.575 -57.145 ;
      RECT 33.475 -53.195 33.575 -53.095 ;
      RECT 33.475 -52.955 33.575 -52.855 ;
      RECT 33.475 -52.715 33.575 -52.615 ;
      RECT 33.475 -52.475 33.575 -52.375 ;
      RECT 33.215 -53.195 33.315 -53.095 ;
      RECT 33.215 -52.955 33.315 -52.855 ;
      RECT 33.215 -52.715 33.315 -52.615 ;
      RECT 33.215 -52.475 33.315 -52.375 ;
      RECT 33.215 -48.5 33.315 -48.4 ;
      RECT 33.215 -45.27 33.315 -45.17 ;
      RECT 33.215 -42.04 33.315 -41.94 ;
      RECT 33.215 -38.81 33.315 -38.71 ;
      RECT 33.215 -35.58 33.315 -35.48 ;
      RECT 33.215 -32.35 33.315 -32.25 ;
      RECT 33.215 -29.12 33.315 -29.02 ;
      RECT 33.215 -25.89 33.315 -25.79 ;
      RECT 33.215 -22.66 33.315 -22.56 ;
      RECT 33.215 -19.43 33.315 -19.33 ;
      RECT 33.215 -16.2 33.315 -16.1 ;
      RECT 33.215 -12.97 33.315 -12.87 ;
      RECT 33.215 -9.74 33.315 -9.64 ;
      RECT 33.215 -6.51 33.315 -6.41 ;
      RECT 33.215 -3.28 33.315 -3.18 ;
      RECT 33.215 -0.05 33.315 0.05 ;
      RECT 33.215 2.245 33.315 2.345 ;
      RECT 33.215 2.485 33.315 2.585 ;
      RECT 33.215 2.725 33.315 2.825 ;
      RECT 33.215 2.965 33.315 3.065 ;
      RECT 32.925 -60.485 33.025 -60.385 ;
      RECT 32.925 -60.285 33.025 -60.185 ;
      RECT 32.925 -59.015 33.025 -58.915 ;
      RECT 32.785 -53.195 32.885 -53.095 ;
      RECT 32.785 -52.955 32.885 -52.855 ;
      RECT 32.785 -52.715 32.885 -52.615 ;
      RECT 32.785 -52.475 32.885 -52.375 ;
      RECT 32.785 -48.5 32.885 -48.4 ;
      RECT 32.785 -45.27 32.885 -45.17 ;
      RECT 32.785 -42.04 32.885 -41.94 ;
      RECT 32.785 -38.81 32.885 -38.71 ;
      RECT 32.785 -35.58 32.885 -35.48 ;
      RECT 32.785 -32.35 32.885 -32.25 ;
      RECT 32.785 -29.12 32.885 -29.02 ;
      RECT 32.785 -25.89 32.885 -25.79 ;
      RECT 32.785 -22.66 32.885 -22.56 ;
      RECT 32.785 -19.43 32.885 -19.33 ;
      RECT 32.785 -16.2 32.885 -16.1 ;
      RECT 32.785 -12.97 32.885 -12.87 ;
      RECT 32.785 -9.74 32.885 -9.64 ;
      RECT 32.785 -6.51 32.885 -6.41 ;
      RECT 32.785 -3.28 32.885 -3.18 ;
      RECT 32.785 -0.05 32.885 0.05 ;
      RECT 32.785 2.245 32.885 2.345 ;
      RECT 32.785 2.485 32.885 2.585 ;
      RECT 32.785 2.725 32.885 2.825 ;
      RECT 32.785 2.965 32.885 3.065 ;
      RECT 32.525 -56.965 32.625 -56.865 ;
      RECT 32.525 -53.195 32.625 -53.095 ;
      RECT 32.525 -52.955 32.625 -52.855 ;
      RECT 32.525 -52.715 32.625 -52.615 ;
      RECT 32.525 -52.475 32.625 -52.375 ;
      RECT 32.335 -60.265 32.435 -60.165 ;
      RECT 32.335 -60.005 32.435 -59.905 ;
      RECT 32.335 -59.03 32.435 -58.93 ;
      RECT 32.335 -58.83 32.435 -58.73 ;
      RECT 32.275 -57.245 32.375 -57.145 ;
      RECT 32.275 -53.195 32.375 -53.095 ;
      RECT 32.275 -52.955 32.375 -52.855 ;
      RECT 32.275 -52.715 32.375 -52.615 ;
      RECT 32.275 -52.475 32.375 -52.375 ;
      RECT 32.035 -57.47 32.135 -57.37 ;
      RECT 32.035 -56.965 32.135 -56.865 ;
      RECT 32.015 -53.195 32.115 -53.095 ;
      RECT 32.015 -52.955 32.115 -52.855 ;
      RECT 32.015 -52.715 32.115 -52.615 ;
      RECT 32.015 -52.475 32.115 -52.375 ;
      RECT 32.015 -48.5 32.115 -48.4 ;
      RECT 32.015 -45.27 32.115 -45.17 ;
      RECT 32.015 -42.04 32.115 -41.94 ;
      RECT 32.015 -38.81 32.115 -38.71 ;
      RECT 32.015 -35.58 32.115 -35.48 ;
      RECT 32.015 -32.35 32.115 -32.25 ;
      RECT 32.015 -29.12 32.115 -29.02 ;
      RECT 32.015 -25.89 32.115 -25.79 ;
      RECT 32.015 -22.66 32.115 -22.56 ;
      RECT 32.015 -19.43 32.115 -19.33 ;
      RECT 32.015 -16.2 32.115 -16.1 ;
      RECT 32.015 -12.97 32.115 -12.87 ;
      RECT 32.015 -9.74 32.115 -9.64 ;
      RECT 32.015 -6.51 32.115 -6.41 ;
      RECT 32.015 -3.28 32.115 -3.18 ;
      RECT 32.015 -0.05 32.115 0.05 ;
      RECT 32.015 2.245 32.115 2.345 ;
      RECT 32.015 2.485 32.115 2.585 ;
      RECT 32.015 2.725 32.115 2.825 ;
      RECT 32.015 2.965 32.115 3.065 ;
      RECT 31.765 -57.875 31.865 -57.775 ;
      RECT 31.585 -53.195 31.685 -53.095 ;
      RECT 31.585 -52.955 31.685 -52.855 ;
      RECT 31.585 -52.715 31.685 -52.615 ;
      RECT 31.585 -52.475 31.685 -52.375 ;
      RECT 31.585 -48.5 31.685 -48.4 ;
      RECT 31.585 -45.27 31.685 -45.17 ;
      RECT 31.585 -42.04 31.685 -41.94 ;
      RECT 31.585 -38.81 31.685 -38.71 ;
      RECT 31.585 -35.58 31.685 -35.48 ;
      RECT 31.585 -32.35 31.685 -32.25 ;
      RECT 31.585 -29.12 31.685 -29.02 ;
      RECT 31.585 -25.89 31.685 -25.79 ;
      RECT 31.585 -22.66 31.685 -22.56 ;
      RECT 31.585 -19.43 31.685 -19.33 ;
      RECT 31.585 -16.2 31.685 -16.1 ;
      RECT 31.585 -12.97 31.685 -12.87 ;
      RECT 31.585 -9.74 31.685 -9.64 ;
      RECT 31.585 -6.51 31.685 -6.41 ;
      RECT 31.585 -3.28 31.685 -3.18 ;
      RECT 31.585 -0.05 31.685 0.05 ;
      RECT 31.585 2.245 31.685 2.345 ;
      RECT 31.585 2.485 31.685 2.585 ;
      RECT 31.585 2.725 31.685 2.825 ;
      RECT 31.585 2.965 31.685 3.065 ;
      RECT 31.44 -57.875 31.54 -57.775 ;
      RECT 31.325 -56.965 31.425 -56.865 ;
      RECT 31.325 -53.195 31.425 -53.095 ;
      RECT 31.325 -52.955 31.425 -52.855 ;
      RECT 31.325 -52.715 31.425 -52.615 ;
      RECT 31.325 -52.475 31.425 -52.375 ;
      RECT 31.075 -57.245 31.175 -57.145 ;
      RECT 31.075 -56.425 31.175 -56.325 ;
      RECT 31.075 -56.185 31.175 -56.085 ;
      RECT 31.075 -55.945 31.175 -55.845 ;
      RECT 31.075 -55.705 31.175 -55.605 ;
      RECT 30.905 -60.485 31.005 -60.385 ;
      RECT 30.905 -60.285 31.005 -60.185 ;
      RECT 30.905 -59.015 31.005 -58.915 ;
      RECT 30.815 -56.425 30.915 -56.325 ;
      RECT 30.815 -56.185 30.915 -56.085 ;
      RECT 30.815 -55.945 30.915 -55.845 ;
      RECT 30.815 -55.705 30.915 -55.605 ;
      RECT 30.815 -48.5 30.915 -48.4 ;
      RECT 30.815 -45.27 30.915 -45.17 ;
      RECT 30.815 -42.04 30.915 -41.94 ;
      RECT 30.815 -38.81 30.915 -38.71 ;
      RECT 30.815 -35.58 30.915 -35.48 ;
      RECT 30.815 -32.35 30.915 -32.25 ;
      RECT 30.815 -29.12 30.915 -29.02 ;
      RECT 30.815 -25.89 30.915 -25.79 ;
      RECT 30.815 -22.66 30.915 -22.56 ;
      RECT 30.815 -19.43 30.915 -19.33 ;
      RECT 30.815 -16.2 30.915 -16.1 ;
      RECT 30.815 -12.97 30.915 -12.87 ;
      RECT 30.815 -9.74 30.915 -9.64 ;
      RECT 30.815 -6.51 30.915 -6.41 ;
      RECT 30.815 -3.28 30.915 -3.18 ;
      RECT 30.815 -0.05 30.915 0.05 ;
      RECT 30.815 2.245 30.915 2.345 ;
      RECT 30.815 2.485 30.915 2.585 ;
      RECT 30.815 2.725 30.915 2.825 ;
      RECT 30.815 2.965 30.915 3.065 ;
      RECT 30.385 -56.425 30.485 -56.325 ;
      RECT 30.385 -56.185 30.485 -56.085 ;
      RECT 30.385 -55.945 30.485 -55.845 ;
      RECT 30.385 -55.705 30.485 -55.605 ;
      RECT 30.385 -48.5 30.485 -48.4 ;
      RECT 30.385 -45.27 30.485 -45.17 ;
      RECT 30.385 -42.04 30.485 -41.94 ;
      RECT 30.385 -38.81 30.485 -38.71 ;
      RECT 30.385 -35.58 30.485 -35.48 ;
      RECT 30.385 -32.35 30.485 -32.25 ;
      RECT 30.385 -29.12 30.485 -29.02 ;
      RECT 30.385 -25.89 30.485 -25.79 ;
      RECT 30.385 -22.66 30.485 -22.56 ;
      RECT 30.385 -19.43 30.485 -19.33 ;
      RECT 30.385 -16.2 30.485 -16.1 ;
      RECT 30.385 -12.97 30.485 -12.87 ;
      RECT 30.385 -9.74 30.485 -9.64 ;
      RECT 30.385 -6.51 30.485 -6.41 ;
      RECT 30.385 -3.28 30.485 -3.18 ;
      RECT 30.385 -0.05 30.485 0.05 ;
      RECT 30.385 2.245 30.485 2.345 ;
      RECT 30.385 2.485 30.485 2.585 ;
      RECT 30.385 2.725 30.485 2.825 ;
      RECT 30.385 2.965 30.485 3.065 ;
      RECT 30.315 -60.265 30.415 -60.165 ;
      RECT 30.315 -60.005 30.415 -59.905 ;
      RECT 30.315 -59.045 30.415 -58.945 ;
      RECT 30.315 -58.845 30.415 -58.745 ;
      RECT 30.125 -56.965 30.225 -56.865 ;
      RECT 30.125 -56.425 30.225 -56.325 ;
      RECT 30.125 -56.185 30.225 -56.085 ;
      RECT 30.125 -55.945 30.225 -55.845 ;
      RECT 30.125 -55.705 30.225 -55.605 ;
      RECT 29.875 -57.245 29.975 -57.145 ;
      RECT 29.875 -56.425 29.975 -56.325 ;
      RECT 29.875 -56.185 29.975 -56.085 ;
      RECT 29.875 -55.945 29.975 -55.845 ;
      RECT 29.875 -55.705 29.975 -55.605 ;
      RECT 29.615 -56.425 29.715 -56.325 ;
      RECT 29.615 -56.185 29.715 -56.085 ;
      RECT 29.615 -55.945 29.715 -55.845 ;
      RECT 29.615 -55.705 29.715 -55.605 ;
      RECT 29.615 -48.5 29.715 -48.4 ;
      RECT 29.615 -45.27 29.715 -45.17 ;
      RECT 29.615 -42.04 29.715 -41.94 ;
      RECT 29.615 -38.81 29.715 -38.71 ;
      RECT 29.615 -35.58 29.715 -35.48 ;
      RECT 29.615 -32.35 29.715 -32.25 ;
      RECT 29.615 -29.12 29.715 -29.02 ;
      RECT 29.615 -25.89 29.715 -25.79 ;
      RECT 29.615 -22.66 29.715 -22.56 ;
      RECT 29.615 -19.43 29.715 -19.33 ;
      RECT 29.615 -16.2 29.715 -16.1 ;
      RECT 29.615 -12.97 29.715 -12.87 ;
      RECT 29.615 -9.74 29.715 -9.64 ;
      RECT 29.615 -6.51 29.715 -6.41 ;
      RECT 29.615 -3.28 29.715 -3.18 ;
      RECT 29.615 -0.05 29.715 0.05 ;
      RECT 29.615 2.245 29.715 2.345 ;
      RECT 29.615 2.485 29.715 2.585 ;
      RECT 29.615 2.725 29.715 2.825 ;
      RECT 29.615 2.965 29.715 3.065 ;
      RECT 29.515 -61.745 29.615 -61.645 ;
      RECT 29.515 -61.545 29.615 -61.445 ;
      RECT 29.185 -56.425 29.285 -56.325 ;
      RECT 29.185 -56.185 29.285 -56.085 ;
      RECT 29.185 -55.945 29.285 -55.845 ;
      RECT 29.185 -55.705 29.285 -55.605 ;
      RECT 29.185 -48.5 29.285 -48.4 ;
      RECT 29.185 -45.27 29.285 -45.17 ;
      RECT 29.185 -42.04 29.285 -41.94 ;
      RECT 29.185 -38.81 29.285 -38.71 ;
      RECT 29.185 -35.58 29.285 -35.48 ;
      RECT 29.185 -32.35 29.285 -32.25 ;
      RECT 29.185 -29.12 29.285 -29.02 ;
      RECT 29.185 -25.89 29.285 -25.79 ;
      RECT 29.185 -22.66 29.285 -22.56 ;
      RECT 29.185 -19.43 29.285 -19.33 ;
      RECT 29.185 -16.2 29.285 -16.1 ;
      RECT 29.185 -12.97 29.285 -12.87 ;
      RECT 29.185 -9.74 29.285 -9.64 ;
      RECT 29.185 -6.51 29.285 -6.41 ;
      RECT 29.185 -3.28 29.285 -3.18 ;
      RECT 29.185 -0.05 29.285 0.05 ;
      RECT 29.185 2.245 29.285 2.345 ;
      RECT 29.185 2.485 29.285 2.585 ;
      RECT 29.185 2.725 29.285 2.825 ;
      RECT 29.185 2.965 29.285 3.065 ;
      RECT 29.165 -60.265 29.265 -60.165 ;
      RECT 29.165 -59.815 29.265 -59.715 ;
      RECT 29.165 -59.015 29.265 -58.915 ;
      RECT 28.925 -61.745 29.025 -61.645 ;
      RECT 28.925 -61.545 29.025 -61.445 ;
      RECT 28.925 -56.965 29.025 -56.865 ;
      RECT 28.925 -56.425 29.025 -56.325 ;
      RECT 28.925 -56.185 29.025 -56.085 ;
      RECT 28.925 -55.945 29.025 -55.845 ;
      RECT 28.925 -55.705 29.025 -55.605 ;
      RECT 28.675 -57.245 28.775 -57.145 ;
      RECT 28.675 -53.195 28.775 -53.095 ;
      RECT 28.675 -52.955 28.775 -52.855 ;
      RECT 28.675 -52.715 28.775 -52.615 ;
      RECT 28.675 -52.475 28.775 -52.375 ;
      RECT 28.415 -53.195 28.515 -53.095 ;
      RECT 28.415 -52.955 28.515 -52.855 ;
      RECT 28.415 -52.715 28.515 -52.615 ;
      RECT 28.415 -52.475 28.515 -52.375 ;
      RECT 28.415 -48.5 28.515 -48.4 ;
      RECT 28.415 -45.27 28.515 -45.17 ;
      RECT 28.415 -42.04 28.515 -41.94 ;
      RECT 28.415 -38.81 28.515 -38.71 ;
      RECT 28.415 -35.58 28.515 -35.48 ;
      RECT 28.415 -32.35 28.515 -32.25 ;
      RECT 28.415 -29.12 28.515 -29.02 ;
      RECT 28.415 -25.89 28.515 -25.79 ;
      RECT 28.415 -22.66 28.515 -22.56 ;
      RECT 28.415 -19.43 28.515 -19.33 ;
      RECT 28.415 -16.2 28.515 -16.1 ;
      RECT 28.415 -12.97 28.515 -12.87 ;
      RECT 28.415 -9.74 28.515 -9.64 ;
      RECT 28.415 -6.51 28.515 -6.41 ;
      RECT 28.415 -3.28 28.515 -3.18 ;
      RECT 28.415 -0.05 28.515 0.05 ;
      RECT 28.415 2.245 28.515 2.345 ;
      RECT 28.415 2.485 28.515 2.585 ;
      RECT 28.415 2.725 28.515 2.825 ;
      RECT 28.415 2.965 28.515 3.065 ;
      RECT 28.125 -60.485 28.225 -60.385 ;
      RECT 28.125 -60.285 28.225 -60.185 ;
      RECT 28.125 -59.015 28.225 -58.915 ;
      RECT 27.985 -53.195 28.085 -53.095 ;
      RECT 27.985 -52.955 28.085 -52.855 ;
      RECT 27.985 -52.715 28.085 -52.615 ;
      RECT 27.985 -52.475 28.085 -52.375 ;
      RECT 27.985 -48.5 28.085 -48.4 ;
      RECT 27.985 -45.27 28.085 -45.17 ;
      RECT 27.985 -42.04 28.085 -41.94 ;
      RECT 27.985 -38.81 28.085 -38.71 ;
      RECT 27.985 -35.58 28.085 -35.48 ;
      RECT 27.985 -32.35 28.085 -32.25 ;
      RECT 27.985 -29.12 28.085 -29.02 ;
      RECT 27.985 -25.89 28.085 -25.79 ;
      RECT 27.985 -22.66 28.085 -22.56 ;
      RECT 27.985 -19.43 28.085 -19.33 ;
      RECT 27.985 -16.2 28.085 -16.1 ;
      RECT 27.985 -12.97 28.085 -12.87 ;
      RECT 27.985 -9.74 28.085 -9.64 ;
      RECT 27.985 -6.51 28.085 -6.41 ;
      RECT 27.985 -3.28 28.085 -3.18 ;
      RECT 27.985 -0.05 28.085 0.05 ;
      RECT 27.985 2.245 28.085 2.345 ;
      RECT 27.985 2.485 28.085 2.585 ;
      RECT 27.985 2.725 28.085 2.825 ;
      RECT 27.985 2.965 28.085 3.065 ;
      RECT 27.725 -56.965 27.825 -56.865 ;
      RECT 27.725 -53.195 27.825 -53.095 ;
      RECT 27.725 -52.955 27.825 -52.855 ;
      RECT 27.725 -52.715 27.825 -52.615 ;
      RECT 27.725 -52.475 27.825 -52.375 ;
      RECT 27.535 -60.265 27.635 -60.165 ;
      RECT 27.535 -60.005 27.635 -59.905 ;
      RECT 27.535 -59.03 27.635 -58.93 ;
      RECT 27.535 -58.83 27.635 -58.73 ;
      RECT 27.475 -57.245 27.575 -57.145 ;
      RECT 27.475 -53.195 27.575 -53.095 ;
      RECT 27.475 -52.955 27.575 -52.855 ;
      RECT 27.475 -52.715 27.575 -52.615 ;
      RECT 27.475 -52.475 27.575 -52.375 ;
      RECT 27.235 -57.47 27.335 -57.37 ;
      RECT 27.235 -56.965 27.335 -56.865 ;
      RECT 27.215 -53.195 27.315 -53.095 ;
      RECT 27.215 -52.955 27.315 -52.855 ;
      RECT 27.215 -52.715 27.315 -52.615 ;
      RECT 27.215 -52.475 27.315 -52.375 ;
      RECT 27.215 -48.5 27.315 -48.4 ;
      RECT 27.215 -45.27 27.315 -45.17 ;
      RECT 27.215 -42.04 27.315 -41.94 ;
      RECT 27.215 -38.81 27.315 -38.71 ;
      RECT 27.215 -35.58 27.315 -35.48 ;
      RECT 27.215 -32.35 27.315 -32.25 ;
      RECT 27.215 -29.12 27.315 -29.02 ;
      RECT 27.215 -25.89 27.315 -25.79 ;
      RECT 27.215 -22.66 27.315 -22.56 ;
      RECT 27.215 -19.43 27.315 -19.33 ;
      RECT 27.215 -16.2 27.315 -16.1 ;
      RECT 27.215 -12.97 27.315 -12.87 ;
      RECT 27.215 -9.74 27.315 -9.64 ;
      RECT 27.215 -6.51 27.315 -6.41 ;
      RECT 27.215 -3.28 27.315 -3.18 ;
      RECT 27.215 -0.05 27.315 0.05 ;
      RECT 27.215 2.245 27.315 2.345 ;
      RECT 27.215 2.485 27.315 2.585 ;
      RECT 27.215 2.725 27.315 2.825 ;
      RECT 27.215 2.965 27.315 3.065 ;
      RECT 26.965 -57.875 27.065 -57.775 ;
      RECT 26.785 -53.195 26.885 -53.095 ;
      RECT 26.785 -52.955 26.885 -52.855 ;
      RECT 26.785 -52.715 26.885 -52.615 ;
      RECT 26.785 -52.475 26.885 -52.375 ;
      RECT 26.785 -48.5 26.885 -48.4 ;
      RECT 26.785 -45.27 26.885 -45.17 ;
      RECT 26.785 -42.04 26.885 -41.94 ;
      RECT 26.785 -38.81 26.885 -38.71 ;
      RECT 26.785 -35.58 26.885 -35.48 ;
      RECT 26.785 -32.35 26.885 -32.25 ;
      RECT 26.785 -29.12 26.885 -29.02 ;
      RECT 26.785 -25.89 26.885 -25.79 ;
      RECT 26.785 -22.66 26.885 -22.56 ;
      RECT 26.785 -19.43 26.885 -19.33 ;
      RECT 26.785 -16.2 26.885 -16.1 ;
      RECT 26.785 -12.97 26.885 -12.87 ;
      RECT 26.785 -9.74 26.885 -9.64 ;
      RECT 26.785 -6.51 26.885 -6.41 ;
      RECT 26.785 -3.28 26.885 -3.18 ;
      RECT 26.785 -0.05 26.885 0.05 ;
      RECT 26.785 2.245 26.885 2.345 ;
      RECT 26.785 2.485 26.885 2.585 ;
      RECT 26.785 2.725 26.885 2.825 ;
      RECT 26.785 2.965 26.885 3.065 ;
      RECT 26.64 -57.875 26.74 -57.775 ;
      RECT 26.525 -56.965 26.625 -56.865 ;
      RECT 26.525 -53.195 26.625 -53.095 ;
      RECT 26.525 -52.955 26.625 -52.855 ;
      RECT 26.525 -52.715 26.625 -52.615 ;
      RECT 26.525 -52.475 26.625 -52.375 ;
      RECT 26.275 -57.245 26.375 -57.145 ;
      RECT 26.275 -56.425 26.375 -56.325 ;
      RECT 26.275 -56.185 26.375 -56.085 ;
      RECT 26.275 -55.945 26.375 -55.845 ;
      RECT 26.275 -55.705 26.375 -55.605 ;
      RECT 26.105 -60.485 26.205 -60.385 ;
      RECT 26.105 -60.285 26.205 -60.185 ;
      RECT 26.105 -59.015 26.205 -58.915 ;
      RECT 26.015 -56.425 26.115 -56.325 ;
      RECT 26.015 -56.185 26.115 -56.085 ;
      RECT 26.015 -55.945 26.115 -55.845 ;
      RECT 26.015 -55.705 26.115 -55.605 ;
      RECT 26.015 -48.5 26.115 -48.4 ;
      RECT 26.015 -45.27 26.115 -45.17 ;
      RECT 26.015 -42.04 26.115 -41.94 ;
      RECT 26.015 -38.81 26.115 -38.71 ;
      RECT 26.015 -35.58 26.115 -35.48 ;
      RECT 26.015 -32.35 26.115 -32.25 ;
      RECT 26.015 -29.12 26.115 -29.02 ;
      RECT 26.015 -25.89 26.115 -25.79 ;
      RECT 26.015 -22.66 26.115 -22.56 ;
      RECT 26.015 -19.43 26.115 -19.33 ;
      RECT 26.015 -16.2 26.115 -16.1 ;
      RECT 26.015 -12.97 26.115 -12.87 ;
      RECT 26.015 -9.74 26.115 -9.64 ;
      RECT 26.015 -6.51 26.115 -6.41 ;
      RECT 26.015 -3.28 26.115 -3.18 ;
      RECT 26.015 -0.05 26.115 0.05 ;
      RECT 26.015 2.245 26.115 2.345 ;
      RECT 26.015 2.485 26.115 2.585 ;
      RECT 26.015 2.725 26.115 2.825 ;
      RECT 26.015 2.965 26.115 3.065 ;
      RECT 25.585 -56.425 25.685 -56.325 ;
      RECT 25.585 -56.185 25.685 -56.085 ;
      RECT 25.585 -55.945 25.685 -55.845 ;
      RECT 25.585 -55.705 25.685 -55.605 ;
      RECT 25.585 -48.5 25.685 -48.4 ;
      RECT 25.585 -45.27 25.685 -45.17 ;
      RECT 25.585 -42.04 25.685 -41.94 ;
      RECT 25.585 -38.81 25.685 -38.71 ;
      RECT 25.585 -35.58 25.685 -35.48 ;
      RECT 25.585 -32.35 25.685 -32.25 ;
      RECT 25.585 -29.12 25.685 -29.02 ;
      RECT 25.585 -25.89 25.685 -25.79 ;
      RECT 25.585 -22.66 25.685 -22.56 ;
      RECT 25.585 -19.43 25.685 -19.33 ;
      RECT 25.585 -16.2 25.685 -16.1 ;
      RECT 25.585 -12.97 25.685 -12.87 ;
      RECT 25.585 -9.74 25.685 -9.64 ;
      RECT 25.585 -6.51 25.685 -6.41 ;
      RECT 25.585 -3.28 25.685 -3.18 ;
      RECT 25.585 -0.05 25.685 0.05 ;
      RECT 25.585 2.245 25.685 2.345 ;
      RECT 25.585 2.485 25.685 2.585 ;
      RECT 25.585 2.725 25.685 2.825 ;
      RECT 25.585 2.965 25.685 3.065 ;
      RECT 25.515 -60.265 25.615 -60.165 ;
      RECT 25.515 -60.005 25.615 -59.905 ;
      RECT 25.515 -59.045 25.615 -58.945 ;
      RECT 25.515 -58.845 25.615 -58.745 ;
      RECT 25.325 -56.965 25.425 -56.865 ;
      RECT 25.325 -56.425 25.425 -56.325 ;
      RECT 25.325 -56.185 25.425 -56.085 ;
      RECT 25.325 -55.945 25.425 -55.845 ;
      RECT 25.325 -55.705 25.425 -55.605 ;
      RECT 25.075 -57.245 25.175 -57.145 ;
      RECT 25.075 -56.425 25.175 -56.325 ;
      RECT 25.075 -56.185 25.175 -56.085 ;
      RECT 25.075 -55.945 25.175 -55.845 ;
      RECT 25.075 -55.705 25.175 -55.605 ;
      RECT 24.815 -56.425 24.915 -56.325 ;
      RECT 24.815 -56.185 24.915 -56.085 ;
      RECT 24.815 -55.945 24.915 -55.845 ;
      RECT 24.815 -55.705 24.915 -55.605 ;
      RECT 24.815 -48.5 24.915 -48.4 ;
      RECT 24.815 -45.27 24.915 -45.17 ;
      RECT 24.815 -42.04 24.915 -41.94 ;
      RECT 24.815 -38.81 24.915 -38.71 ;
      RECT 24.815 -35.58 24.915 -35.48 ;
      RECT 24.815 -32.35 24.915 -32.25 ;
      RECT 24.815 -29.12 24.915 -29.02 ;
      RECT 24.815 -25.89 24.915 -25.79 ;
      RECT 24.815 -22.66 24.915 -22.56 ;
      RECT 24.815 -19.43 24.915 -19.33 ;
      RECT 24.815 -16.2 24.915 -16.1 ;
      RECT 24.815 -12.97 24.915 -12.87 ;
      RECT 24.815 -9.74 24.915 -9.64 ;
      RECT 24.815 -6.51 24.915 -6.41 ;
      RECT 24.815 -3.28 24.915 -3.18 ;
      RECT 24.815 -0.05 24.915 0.05 ;
      RECT 24.815 2.245 24.915 2.345 ;
      RECT 24.815 2.485 24.915 2.585 ;
      RECT 24.815 2.725 24.915 2.825 ;
      RECT 24.815 2.965 24.915 3.065 ;
      RECT 24.715 -61.745 24.815 -61.645 ;
      RECT 24.715 -61.545 24.815 -61.445 ;
      RECT 24.385 -56.425 24.485 -56.325 ;
      RECT 24.385 -56.185 24.485 -56.085 ;
      RECT 24.385 -55.945 24.485 -55.845 ;
      RECT 24.385 -55.705 24.485 -55.605 ;
      RECT 24.385 -48.5 24.485 -48.4 ;
      RECT 24.385 -45.27 24.485 -45.17 ;
      RECT 24.385 -42.04 24.485 -41.94 ;
      RECT 24.385 -38.81 24.485 -38.71 ;
      RECT 24.385 -35.58 24.485 -35.48 ;
      RECT 24.385 -32.35 24.485 -32.25 ;
      RECT 24.385 -29.12 24.485 -29.02 ;
      RECT 24.385 -25.89 24.485 -25.79 ;
      RECT 24.385 -22.66 24.485 -22.56 ;
      RECT 24.385 -19.43 24.485 -19.33 ;
      RECT 24.385 -16.2 24.485 -16.1 ;
      RECT 24.385 -12.97 24.485 -12.87 ;
      RECT 24.385 -9.74 24.485 -9.64 ;
      RECT 24.385 -6.51 24.485 -6.41 ;
      RECT 24.385 -3.28 24.485 -3.18 ;
      RECT 24.385 -0.05 24.485 0.05 ;
      RECT 24.385 2.245 24.485 2.345 ;
      RECT 24.385 2.485 24.485 2.585 ;
      RECT 24.385 2.725 24.485 2.825 ;
      RECT 24.385 2.965 24.485 3.065 ;
      RECT 24.365 -60.265 24.465 -60.165 ;
      RECT 24.365 -59.815 24.465 -59.715 ;
      RECT 24.365 -59.015 24.465 -58.915 ;
      RECT 24.125 -61.745 24.225 -61.645 ;
      RECT 24.125 -61.545 24.225 -61.445 ;
      RECT 24.125 -56.965 24.225 -56.865 ;
      RECT 24.125 -56.425 24.225 -56.325 ;
      RECT 24.125 -56.185 24.225 -56.085 ;
      RECT 24.125 -55.945 24.225 -55.845 ;
      RECT 24.125 -55.705 24.225 -55.605 ;
      RECT 23.875 -57.245 23.975 -57.145 ;
      RECT 23.875 -53.195 23.975 -53.095 ;
      RECT 23.875 -52.955 23.975 -52.855 ;
      RECT 23.875 -52.715 23.975 -52.615 ;
      RECT 23.875 -52.475 23.975 -52.375 ;
      RECT 23.615 -53.195 23.715 -53.095 ;
      RECT 23.615 -52.955 23.715 -52.855 ;
      RECT 23.615 -52.715 23.715 -52.615 ;
      RECT 23.615 -52.475 23.715 -52.375 ;
      RECT 23.615 -48.5 23.715 -48.4 ;
      RECT 23.615 -45.27 23.715 -45.17 ;
      RECT 23.615 -42.04 23.715 -41.94 ;
      RECT 23.615 -38.81 23.715 -38.71 ;
      RECT 23.615 -35.58 23.715 -35.48 ;
      RECT 23.615 -32.35 23.715 -32.25 ;
      RECT 23.615 -29.12 23.715 -29.02 ;
      RECT 23.615 -25.89 23.715 -25.79 ;
      RECT 23.615 -22.66 23.715 -22.56 ;
      RECT 23.615 -19.43 23.715 -19.33 ;
      RECT 23.615 -16.2 23.715 -16.1 ;
      RECT 23.615 -12.97 23.715 -12.87 ;
      RECT 23.615 -9.74 23.715 -9.64 ;
      RECT 23.615 -6.51 23.715 -6.41 ;
      RECT 23.615 -3.28 23.715 -3.18 ;
      RECT 23.615 -0.05 23.715 0.05 ;
      RECT 23.615 2.245 23.715 2.345 ;
      RECT 23.615 2.485 23.715 2.585 ;
      RECT 23.615 2.725 23.715 2.825 ;
      RECT 23.615 2.965 23.715 3.065 ;
      RECT 23.325 -60.485 23.425 -60.385 ;
      RECT 23.325 -60.285 23.425 -60.185 ;
      RECT 23.325 -59.015 23.425 -58.915 ;
      RECT 23.185 -53.195 23.285 -53.095 ;
      RECT 23.185 -52.955 23.285 -52.855 ;
      RECT 23.185 -52.715 23.285 -52.615 ;
      RECT 23.185 -52.475 23.285 -52.375 ;
      RECT 23.185 -48.5 23.285 -48.4 ;
      RECT 23.185 -45.27 23.285 -45.17 ;
      RECT 23.185 -42.04 23.285 -41.94 ;
      RECT 23.185 -38.81 23.285 -38.71 ;
      RECT 23.185 -35.58 23.285 -35.48 ;
      RECT 23.185 -32.35 23.285 -32.25 ;
      RECT 23.185 -29.12 23.285 -29.02 ;
      RECT 23.185 -25.89 23.285 -25.79 ;
      RECT 23.185 -22.66 23.285 -22.56 ;
      RECT 23.185 -19.43 23.285 -19.33 ;
      RECT 23.185 -16.2 23.285 -16.1 ;
      RECT 23.185 -12.97 23.285 -12.87 ;
      RECT 23.185 -9.74 23.285 -9.64 ;
      RECT 23.185 -6.51 23.285 -6.41 ;
      RECT 23.185 -3.28 23.285 -3.18 ;
      RECT 23.185 -0.05 23.285 0.05 ;
      RECT 23.185 2.245 23.285 2.345 ;
      RECT 23.185 2.485 23.285 2.585 ;
      RECT 23.185 2.725 23.285 2.825 ;
      RECT 23.185 2.965 23.285 3.065 ;
      RECT 22.925 -56.965 23.025 -56.865 ;
      RECT 22.925 -53.195 23.025 -53.095 ;
      RECT 22.925 -52.955 23.025 -52.855 ;
      RECT 22.925 -52.715 23.025 -52.615 ;
      RECT 22.925 -52.475 23.025 -52.375 ;
      RECT 22.735 -60.265 22.835 -60.165 ;
      RECT 22.735 -60.005 22.835 -59.905 ;
      RECT 22.735 -59.03 22.835 -58.93 ;
      RECT 22.735 -58.83 22.835 -58.73 ;
      RECT 22.675 -57.245 22.775 -57.145 ;
      RECT 22.675 -53.195 22.775 -53.095 ;
      RECT 22.675 -52.955 22.775 -52.855 ;
      RECT 22.675 -52.715 22.775 -52.615 ;
      RECT 22.675 -52.475 22.775 -52.375 ;
      RECT 22.435 -57.47 22.535 -57.37 ;
      RECT 22.435 -56.965 22.535 -56.865 ;
      RECT 22.415 -53.195 22.515 -53.095 ;
      RECT 22.415 -52.955 22.515 -52.855 ;
      RECT 22.415 -52.715 22.515 -52.615 ;
      RECT 22.415 -52.475 22.515 -52.375 ;
      RECT 22.415 -48.5 22.515 -48.4 ;
      RECT 22.415 -45.27 22.515 -45.17 ;
      RECT 22.415 -42.04 22.515 -41.94 ;
      RECT 22.415 -38.81 22.515 -38.71 ;
      RECT 22.415 -35.58 22.515 -35.48 ;
      RECT 22.415 -32.35 22.515 -32.25 ;
      RECT 22.415 -29.12 22.515 -29.02 ;
      RECT 22.415 -25.89 22.515 -25.79 ;
      RECT 22.415 -22.66 22.515 -22.56 ;
      RECT 22.415 -19.43 22.515 -19.33 ;
      RECT 22.415 -16.2 22.515 -16.1 ;
      RECT 22.415 -12.97 22.515 -12.87 ;
      RECT 22.415 -9.74 22.515 -9.64 ;
      RECT 22.415 -6.51 22.515 -6.41 ;
      RECT 22.415 -3.28 22.515 -3.18 ;
      RECT 22.415 -0.05 22.515 0.05 ;
      RECT 22.415 2.245 22.515 2.345 ;
      RECT 22.415 2.485 22.515 2.585 ;
      RECT 22.415 2.725 22.515 2.825 ;
      RECT 22.415 2.965 22.515 3.065 ;
      RECT 22.165 -57.875 22.265 -57.775 ;
      RECT 21.985 -53.195 22.085 -53.095 ;
      RECT 21.985 -52.955 22.085 -52.855 ;
      RECT 21.985 -52.715 22.085 -52.615 ;
      RECT 21.985 -52.475 22.085 -52.375 ;
      RECT 21.985 -48.5 22.085 -48.4 ;
      RECT 21.985 -45.27 22.085 -45.17 ;
      RECT 21.985 -42.04 22.085 -41.94 ;
      RECT 21.985 -38.81 22.085 -38.71 ;
      RECT 21.985 -35.58 22.085 -35.48 ;
      RECT 21.985 -32.35 22.085 -32.25 ;
      RECT 21.985 -29.12 22.085 -29.02 ;
      RECT 21.985 -25.89 22.085 -25.79 ;
      RECT 21.985 -22.66 22.085 -22.56 ;
      RECT 21.985 -19.43 22.085 -19.33 ;
      RECT 21.985 -16.2 22.085 -16.1 ;
      RECT 21.985 -12.97 22.085 -12.87 ;
      RECT 21.985 -9.74 22.085 -9.64 ;
      RECT 21.985 -6.51 22.085 -6.41 ;
      RECT 21.985 -3.28 22.085 -3.18 ;
      RECT 21.985 -0.05 22.085 0.05 ;
      RECT 21.985 2.245 22.085 2.345 ;
      RECT 21.985 2.485 22.085 2.585 ;
      RECT 21.985 2.725 22.085 2.825 ;
      RECT 21.985 2.965 22.085 3.065 ;
      RECT 21.84 -57.875 21.94 -57.775 ;
      RECT 21.725 -56.965 21.825 -56.865 ;
      RECT 21.725 -53.195 21.825 -53.095 ;
      RECT 21.725 -52.955 21.825 -52.855 ;
      RECT 21.725 -52.715 21.825 -52.615 ;
      RECT 21.725 -52.475 21.825 -52.375 ;
      RECT 21.475 -57.245 21.575 -57.145 ;
      RECT 21.475 -56.425 21.575 -56.325 ;
      RECT 21.475 -56.185 21.575 -56.085 ;
      RECT 21.475 -55.945 21.575 -55.845 ;
      RECT 21.475 -55.705 21.575 -55.605 ;
      RECT 21.305 -60.485 21.405 -60.385 ;
      RECT 21.305 -60.285 21.405 -60.185 ;
      RECT 21.305 -59.015 21.405 -58.915 ;
      RECT 21.215 -56.425 21.315 -56.325 ;
      RECT 21.215 -56.185 21.315 -56.085 ;
      RECT 21.215 -55.945 21.315 -55.845 ;
      RECT 21.215 -55.705 21.315 -55.605 ;
      RECT 21.215 -48.5 21.315 -48.4 ;
      RECT 21.215 -45.27 21.315 -45.17 ;
      RECT 21.215 -42.04 21.315 -41.94 ;
      RECT 21.215 -38.81 21.315 -38.71 ;
      RECT 21.215 -35.58 21.315 -35.48 ;
      RECT 21.215 -32.35 21.315 -32.25 ;
      RECT 21.215 -29.12 21.315 -29.02 ;
      RECT 21.215 -25.89 21.315 -25.79 ;
      RECT 21.215 -22.66 21.315 -22.56 ;
      RECT 21.215 -19.43 21.315 -19.33 ;
      RECT 21.215 -16.2 21.315 -16.1 ;
      RECT 21.215 -12.97 21.315 -12.87 ;
      RECT 21.215 -9.74 21.315 -9.64 ;
      RECT 21.215 -6.51 21.315 -6.41 ;
      RECT 21.215 -3.28 21.315 -3.18 ;
      RECT 21.215 -0.05 21.315 0.05 ;
      RECT 21.215 2.245 21.315 2.345 ;
      RECT 21.215 2.485 21.315 2.585 ;
      RECT 21.215 2.725 21.315 2.825 ;
      RECT 21.215 2.965 21.315 3.065 ;
      RECT 20.785 -56.425 20.885 -56.325 ;
      RECT 20.785 -56.185 20.885 -56.085 ;
      RECT 20.785 -55.945 20.885 -55.845 ;
      RECT 20.785 -55.705 20.885 -55.605 ;
      RECT 20.785 -48.5 20.885 -48.4 ;
      RECT 20.785 -45.27 20.885 -45.17 ;
      RECT 20.785 -42.04 20.885 -41.94 ;
      RECT 20.785 -38.81 20.885 -38.71 ;
      RECT 20.785 -35.58 20.885 -35.48 ;
      RECT 20.785 -32.35 20.885 -32.25 ;
      RECT 20.785 -29.12 20.885 -29.02 ;
      RECT 20.785 -25.89 20.885 -25.79 ;
      RECT 20.785 -22.66 20.885 -22.56 ;
      RECT 20.785 -19.43 20.885 -19.33 ;
      RECT 20.785 -16.2 20.885 -16.1 ;
      RECT 20.785 -12.97 20.885 -12.87 ;
      RECT 20.785 -9.74 20.885 -9.64 ;
      RECT 20.785 -6.51 20.885 -6.41 ;
      RECT 20.785 -3.28 20.885 -3.18 ;
      RECT 20.785 -0.05 20.885 0.05 ;
      RECT 20.785 2.245 20.885 2.345 ;
      RECT 20.785 2.485 20.885 2.585 ;
      RECT 20.785 2.725 20.885 2.825 ;
      RECT 20.785 2.965 20.885 3.065 ;
      RECT 20.715 -60.265 20.815 -60.165 ;
      RECT 20.715 -60.005 20.815 -59.905 ;
      RECT 20.715 -59.045 20.815 -58.945 ;
      RECT 20.715 -58.845 20.815 -58.745 ;
      RECT 20.525 -56.965 20.625 -56.865 ;
      RECT 20.525 -56.425 20.625 -56.325 ;
      RECT 20.525 -56.185 20.625 -56.085 ;
      RECT 20.525 -55.945 20.625 -55.845 ;
      RECT 20.525 -55.705 20.625 -55.605 ;
      RECT 20.275 -57.245 20.375 -57.145 ;
      RECT 20.275 -56.425 20.375 -56.325 ;
      RECT 20.275 -56.185 20.375 -56.085 ;
      RECT 20.275 -55.945 20.375 -55.845 ;
      RECT 20.275 -55.705 20.375 -55.605 ;
      RECT 20.015 -56.425 20.115 -56.325 ;
      RECT 20.015 -56.185 20.115 -56.085 ;
      RECT 20.015 -55.945 20.115 -55.845 ;
      RECT 20.015 -55.705 20.115 -55.605 ;
      RECT 20.015 -48.5 20.115 -48.4 ;
      RECT 20.015 -45.27 20.115 -45.17 ;
      RECT 20.015 -42.04 20.115 -41.94 ;
      RECT 20.015 -38.81 20.115 -38.71 ;
      RECT 20.015 -35.58 20.115 -35.48 ;
      RECT 20.015 -32.35 20.115 -32.25 ;
      RECT 20.015 -29.12 20.115 -29.02 ;
      RECT 20.015 -25.89 20.115 -25.79 ;
      RECT 20.015 -22.66 20.115 -22.56 ;
      RECT 20.015 -19.43 20.115 -19.33 ;
      RECT 20.015 -16.2 20.115 -16.1 ;
      RECT 20.015 -12.97 20.115 -12.87 ;
      RECT 20.015 -9.74 20.115 -9.64 ;
      RECT 20.015 -6.51 20.115 -6.41 ;
      RECT 20.015 -3.28 20.115 -3.18 ;
      RECT 20.015 -0.05 20.115 0.05 ;
      RECT 20.015 2.245 20.115 2.345 ;
      RECT 20.015 2.485 20.115 2.585 ;
      RECT 20.015 2.725 20.115 2.825 ;
      RECT 20.015 2.965 20.115 3.065 ;
      RECT 19.915 -61.745 20.015 -61.645 ;
      RECT 19.915 -61.545 20.015 -61.445 ;
      RECT 19.585 -56.425 19.685 -56.325 ;
      RECT 19.585 -56.185 19.685 -56.085 ;
      RECT 19.585 -55.945 19.685 -55.845 ;
      RECT 19.585 -55.705 19.685 -55.605 ;
      RECT 19.585 -48.5 19.685 -48.4 ;
      RECT 19.585 -45.27 19.685 -45.17 ;
      RECT 19.585 -42.04 19.685 -41.94 ;
      RECT 19.585 -38.81 19.685 -38.71 ;
      RECT 19.585 -35.58 19.685 -35.48 ;
      RECT 19.585 -32.35 19.685 -32.25 ;
      RECT 19.585 -29.12 19.685 -29.02 ;
      RECT 19.585 -25.89 19.685 -25.79 ;
      RECT 19.585 -22.66 19.685 -22.56 ;
      RECT 19.585 -19.43 19.685 -19.33 ;
      RECT 19.585 -16.2 19.685 -16.1 ;
      RECT 19.585 -12.97 19.685 -12.87 ;
      RECT 19.585 -9.74 19.685 -9.64 ;
      RECT 19.585 -6.51 19.685 -6.41 ;
      RECT 19.585 -3.28 19.685 -3.18 ;
      RECT 19.585 -0.05 19.685 0.05 ;
      RECT 19.585 2.245 19.685 2.345 ;
      RECT 19.585 2.485 19.685 2.585 ;
      RECT 19.585 2.725 19.685 2.825 ;
      RECT 19.585 2.965 19.685 3.065 ;
      RECT 19.565 -60.265 19.665 -60.165 ;
      RECT 19.565 -59.815 19.665 -59.715 ;
      RECT 19.565 -59.015 19.665 -58.915 ;
      RECT 19.325 -61.745 19.425 -61.645 ;
      RECT 19.325 -61.545 19.425 -61.445 ;
      RECT 19.325 -56.965 19.425 -56.865 ;
      RECT 19.325 -56.425 19.425 -56.325 ;
      RECT 19.325 -56.185 19.425 -56.085 ;
      RECT 19.325 -55.945 19.425 -55.845 ;
      RECT 19.325 -55.705 19.425 -55.605 ;
      RECT 19.075 -57.245 19.175 -57.145 ;
      RECT 19.075 -53.195 19.175 -53.095 ;
      RECT 19.075 -52.955 19.175 -52.855 ;
      RECT 19.075 -52.715 19.175 -52.615 ;
      RECT 19.075 -52.475 19.175 -52.375 ;
      RECT 18.815 -53.195 18.915 -53.095 ;
      RECT 18.815 -52.955 18.915 -52.855 ;
      RECT 18.815 -52.715 18.915 -52.615 ;
      RECT 18.815 -52.475 18.915 -52.375 ;
      RECT 18.815 -48.5 18.915 -48.4 ;
      RECT 18.815 -45.27 18.915 -45.17 ;
      RECT 18.815 -42.04 18.915 -41.94 ;
      RECT 18.815 -38.81 18.915 -38.71 ;
      RECT 18.815 -35.58 18.915 -35.48 ;
      RECT 18.815 -32.35 18.915 -32.25 ;
      RECT 18.815 -29.12 18.915 -29.02 ;
      RECT 18.815 -25.89 18.915 -25.79 ;
      RECT 18.815 -22.66 18.915 -22.56 ;
      RECT 18.815 -19.43 18.915 -19.33 ;
      RECT 18.815 -16.2 18.915 -16.1 ;
      RECT 18.815 -12.97 18.915 -12.87 ;
      RECT 18.815 -9.74 18.915 -9.64 ;
      RECT 18.815 -6.51 18.915 -6.41 ;
      RECT 18.815 -3.28 18.915 -3.18 ;
      RECT 18.815 -0.05 18.915 0.05 ;
      RECT 18.815 2.245 18.915 2.345 ;
      RECT 18.815 2.485 18.915 2.585 ;
      RECT 18.815 2.725 18.915 2.825 ;
      RECT 18.815 2.965 18.915 3.065 ;
      RECT 18.525 -60.485 18.625 -60.385 ;
      RECT 18.525 -60.285 18.625 -60.185 ;
      RECT 18.525 -59.015 18.625 -58.915 ;
      RECT 18.385 -53.195 18.485 -53.095 ;
      RECT 18.385 -52.955 18.485 -52.855 ;
      RECT 18.385 -52.715 18.485 -52.615 ;
      RECT 18.385 -52.475 18.485 -52.375 ;
      RECT 18.385 -48.5 18.485 -48.4 ;
      RECT 18.385 -45.27 18.485 -45.17 ;
      RECT 18.385 -42.04 18.485 -41.94 ;
      RECT 18.385 -38.81 18.485 -38.71 ;
      RECT 18.385 -35.58 18.485 -35.48 ;
      RECT 18.385 -32.35 18.485 -32.25 ;
      RECT 18.385 -29.12 18.485 -29.02 ;
      RECT 18.385 -25.89 18.485 -25.79 ;
      RECT 18.385 -22.66 18.485 -22.56 ;
      RECT 18.385 -19.43 18.485 -19.33 ;
      RECT 18.385 -16.2 18.485 -16.1 ;
      RECT 18.385 -12.97 18.485 -12.87 ;
      RECT 18.385 -9.74 18.485 -9.64 ;
      RECT 18.385 -6.51 18.485 -6.41 ;
      RECT 18.385 -3.28 18.485 -3.18 ;
      RECT 18.385 -0.05 18.485 0.05 ;
      RECT 18.385 2.245 18.485 2.345 ;
      RECT 18.385 2.485 18.485 2.585 ;
      RECT 18.385 2.725 18.485 2.825 ;
      RECT 18.385 2.965 18.485 3.065 ;
      RECT 18.125 -56.965 18.225 -56.865 ;
      RECT 18.125 -53.195 18.225 -53.095 ;
      RECT 18.125 -52.955 18.225 -52.855 ;
      RECT 18.125 -52.715 18.225 -52.615 ;
      RECT 18.125 -52.475 18.225 -52.375 ;
      RECT 17.935 -60.265 18.035 -60.165 ;
      RECT 17.935 -60.005 18.035 -59.905 ;
      RECT 17.935 -59.03 18.035 -58.93 ;
      RECT 17.935 -58.83 18.035 -58.73 ;
      RECT 17.875 -57.245 17.975 -57.145 ;
      RECT 17.875 -53.195 17.975 -53.095 ;
      RECT 17.875 -52.955 17.975 -52.855 ;
      RECT 17.875 -52.715 17.975 -52.615 ;
      RECT 17.875 -52.475 17.975 -52.375 ;
      RECT 17.635 -57.47 17.735 -57.37 ;
      RECT 17.635 -56.965 17.735 -56.865 ;
      RECT 17.615 -53.195 17.715 -53.095 ;
      RECT 17.615 -52.955 17.715 -52.855 ;
      RECT 17.615 -52.715 17.715 -52.615 ;
      RECT 17.615 -52.475 17.715 -52.375 ;
      RECT 17.615 -48.5 17.715 -48.4 ;
      RECT 17.615 -45.27 17.715 -45.17 ;
      RECT 17.615 -42.04 17.715 -41.94 ;
      RECT 17.615 -38.81 17.715 -38.71 ;
      RECT 17.615 -35.58 17.715 -35.48 ;
      RECT 17.615 -32.35 17.715 -32.25 ;
      RECT 17.615 -29.12 17.715 -29.02 ;
      RECT 17.615 -25.89 17.715 -25.79 ;
      RECT 17.615 -22.66 17.715 -22.56 ;
      RECT 17.615 -19.43 17.715 -19.33 ;
      RECT 17.615 -16.2 17.715 -16.1 ;
      RECT 17.615 -12.97 17.715 -12.87 ;
      RECT 17.615 -9.74 17.715 -9.64 ;
      RECT 17.615 -6.51 17.715 -6.41 ;
      RECT 17.615 -3.28 17.715 -3.18 ;
      RECT 17.615 -0.05 17.715 0.05 ;
      RECT 17.615 2.245 17.715 2.345 ;
      RECT 17.615 2.485 17.715 2.585 ;
      RECT 17.615 2.725 17.715 2.825 ;
      RECT 17.615 2.965 17.715 3.065 ;
      RECT 17.365 -57.875 17.465 -57.775 ;
      RECT 17.185 -53.195 17.285 -53.095 ;
      RECT 17.185 -52.955 17.285 -52.855 ;
      RECT 17.185 -52.715 17.285 -52.615 ;
      RECT 17.185 -52.475 17.285 -52.375 ;
      RECT 17.185 -48.5 17.285 -48.4 ;
      RECT 17.185 -45.27 17.285 -45.17 ;
      RECT 17.185 -42.04 17.285 -41.94 ;
      RECT 17.185 -38.81 17.285 -38.71 ;
      RECT 17.185 -35.58 17.285 -35.48 ;
      RECT 17.185 -32.35 17.285 -32.25 ;
      RECT 17.185 -29.12 17.285 -29.02 ;
      RECT 17.185 -25.89 17.285 -25.79 ;
      RECT 17.185 -22.66 17.285 -22.56 ;
      RECT 17.185 -19.43 17.285 -19.33 ;
      RECT 17.185 -16.2 17.285 -16.1 ;
      RECT 17.185 -12.97 17.285 -12.87 ;
      RECT 17.185 -9.74 17.285 -9.64 ;
      RECT 17.185 -6.51 17.285 -6.41 ;
      RECT 17.185 -3.28 17.285 -3.18 ;
      RECT 17.185 -0.05 17.285 0.05 ;
      RECT 17.185 2.245 17.285 2.345 ;
      RECT 17.185 2.485 17.285 2.585 ;
      RECT 17.185 2.725 17.285 2.825 ;
      RECT 17.185 2.965 17.285 3.065 ;
      RECT 17.04 -57.875 17.14 -57.775 ;
      RECT 16.925 -56.965 17.025 -56.865 ;
      RECT 16.925 -53.195 17.025 -53.095 ;
      RECT 16.925 -52.955 17.025 -52.855 ;
      RECT 16.925 -52.715 17.025 -52.615 ;
      RECT 16.925 -52.475 17.025 -52.375 ;
      RECT 16.675 -57.245 16.775 -57.145 ;
      RECT 16.675 -56.425 16.775 -56.325 ;
      RECT 16.675 -56.185 16.775 -56.085 ;
      RECT 16.675 -55.945 16.775 -55.845 ;
      RECT 16.675 -55.705 16.775 -55.605 ;
      RECT 16.505 -60.485 16.605 -60.385 ;
      RECT 16.505 -60.285 16.605 -60.185 ;
      RECT 16.505 -59.015 16.605 -58.915 ;
      RECT 16.415 -56.425 16.515 -56.325 ;
      RECT 16.415 -56.185 16.515 -56.085 ;
      RECT 16.415 -55.945 16.515 -55.845 ;
      RECT 16.415 -55.705 16.515 -55.605 ;
      RECT 16.415 -48.5 16.515 -48.4 ;
      RECT 16.415 -45.27 16.515 -45.17 ;
      RECT 16.415 -42.04 16.515 -41.94 ;
      RECT 16.415 -38.81 16.515 -38.71 ;
      RECT 16.415 -35.58 16.515 -35.48 ;
      RECT 16.415 -32.35 16.515 -32.25 ;
      RECT 16.415 -29.12 16.515 -29.02 ;
      RECT 16.415 -25.89 16.515 -25.79 ;
      RECT 16.415 -22.66 16.515 -22.56 ;
      RECT 16.415 -19.43 16.515 -19.33 ;
      RECT 16.415 -16.2 16.515 -16.1 ;
      RECT 16.415 -12.97 16.515 -12.87 ;
      RECT 16.415 -9.74 16.515 -9.64 ;
      RECT 16.415 -6.51 16.515 -6.41 ;
      RECT 16.415 -3.28 16.515 -3.18 ;
      RECT 16.415 -0.05 16.515 0.05 ;
      RECT 16.415 2.245 16.515 2.345 ;
      RECT 16.415 2.485 16.515 2.585 ;
      RECT 16.415 2.725 16.515 2.825 ;
      RECT 16.415 2.965 16.515 3.065 ;
      RECT 15.985 -56.425 16.085 -56.325 ;
      RECT 15.985 -56.185 16.085 -56.085 ;
      RECT 15.985 -55.945 16.085 -55.845 ;
      RECT 15.985 -55.705 16.085 -55.605 ;
      RECT 15.985 -48.5 16.085 -48.4 ;
      RECT 15.985 -45.27 16.085 -45.17 ;
      RECT 15.985 -42.04 16.085 -41.94 ;
      RECT 15.985 -38.81 16.085 -38.71 ;
      RECT 15.985 -35.58 16.085 -35.48 ;
      RECT 15.985 -32.35 16.085 -32.25 ;
      RECT 15.985 -29.12 16.085 -29.02 ;
      RECT 15.985 -25.89 16.085 -25.79 ;
      RECT 15.985 -22.66 16.085 -22.56 ;
      RECT 15.985 -19.43 16.085 -19.33 ;
      RECT 15.985 -16.2 16.085 -16.1 ;
      RECT 15.985 -12.97 16.085 -12.87 ;
      RECT 15.985 -9.74 16.085 -9.64 ;
      RECT 15.985 -6.51 16.085 -6.41 ;
      RECT 15.985 -3.28 16.085 -3.18 ;
      RECT 15.985 -0.05 16.085 0.05 ;
      RECT 15.985 2.245 16.085 2.345 ;
      RECT 15.985 2.485 16.085 2.585 ;
      RECT 15.985 2.725 16.085 2.825 ;
      RECT 15.985 2.965 16.085 3.065 ;
      RECT 15.915 -60.265 16.015 -60.165 ;
      RECT 15.915 -60.005 16.015 -59.905 ;
      RECT 15.915 -59.045 16.015 -58.945 ;
      RECT 15.915 -58.845 16.015 -58.745 ;
      RECT 15.725 -56.965 15.825 -56.865 ;
      RECT 15.725 -56.425 15.825 -56.325 ;
      RECT 15.725 -56.185 15.825 -56.085 ;
      RECT 15.725 -55.945 15.825 -55.845 ;
      RECT 15.725 -55.705 15.825 -55.605 ;
      RECT 15.475 -57.245 15.575 -57.145 ;
      RECT 15.475 -56.425 15.575 -56.325 ;
      RECT 15.475 -56.185 15.575 -56.085 ;
      RECT 15.475 -55.945 15.575 -55.845 ;
      RECT 15.475 -55.705 15.575 -55.605 ;
      RECT 15.215 -56.425 15.315 -56.325 ;
      RECT 15.215 -56.185 15.315 -56.085 ;
      RECT 15.215 -55.945 15.315 -55.845 ;
      RECT 15.215 -55.705 15.315 -55.605 ;
      RECT 15.215 -48.5 15.315 -48.4 ;
      RECT 15.215 -45.27 15.315 -45.17 ;
      RECT 15.215 -42.04 15.315 -41.94 ;
      RECT 15.215 -38.81 15.315 -38.71 ;
      RECT 15.215 -35.58 15.315 -35.48 ;
      RECT 15.215 -32.35 15.315 -32.25 ;
      RECT 15.215 -29.12 15.315 -29.02 ;
      RECT 15.215 -25.89 15.315 -25.79 ;
      RECT 15.215 -22.66 15.315 -22.56 ;
      RECT 15.215 -19.43 15.315 -19.33 ;
      RECT 15.215 -16.2 15.315 -16.1 ;
      RECT 15.215 -12.97 15.315 -12.87 ;
      RECT 15.215 -9.74 15.315 -9.64 ;
      RECT 15.215 -6.51 15.315 -6.41 ;
      RECT 15.215 -3.28 15.315 -3.18 ;
      RECT 15.215 -0.05 15.315 0.05 ;
      RECT 15.215 2.245 15.315 2.345 ;
      RECT 15.215 2.485 15.315 2.585 ;
      RECT 15.215 2.725 15.315 2.825 ;
      RECT 15.215 2.965 15.315 3.065 ;
      RECT 15.115 -61.745 15.215 -61.645 ;
      RECT 15.115 -61.545 15.215 -61.445 ;
      RECT 14.785 -56.425 14.885 -56.325 ;
      RECT 14.785 -56.185 14.885 -56.085 ;
      RECT 14.785 -55.945 14.885 -55.845 ;
      RECT 14.785 -55.705 14.885 -55.605 ;
      RECT 14.785 -48.5 14.885 -48.4 ;
      RECT 14.785 -45.27 14.885 -45.17 ;
      RECT 14.785 -42.04 14.885 -41.94 ;
      RECT 14.785 -38.81 14.885 -38.71 ;
      RECT 14.785 -35.58 14.885 -35.48 ;
      RECT 14.785 -32.35 14.885 -32.25 ;
      RECT 14.785 -29.12 14.885 -29.02 ;
      RECT 14.785 -25.89 14.885 -25.79 ;
      RECT 14.785 -22.66 14.885 -22.56 ;
      RECT 14.785 -19.43 14.885 -19.33 ;
      RECT 14.785 -16.2 14.885 -16.1 ;
      RECT 14.785 -12.97 14.885 -12.87 ;
      RECT 14.785 -9.74 14.885 -9.64 ;
      RECT 14.785 -6.51 14.885 -6.41 ;
      RECT 14.785 -3.28 14.885 -3.18 ;
      RECT 14.785 -0.05 14.885 0.05 ;
      RECT 14.785 2.245 14.885 2.345 ;
      RECT 14.785 2.485 14.885 2.585 ;
      RECT 14.785 2.725 14.885 2.825 ;
      RECT 14.785 2.965 14.885 3.065 ;
      RECT 14.765 -60.265 14.865 -60.165 ;
      RECT 14.765 -59.815 14.865 -59.715 ;
      RECT 14.765 -59.015 14.865 -58.915 ;
      RECT 14.525 -61.745 14.625 -61.645 ;
      RECT 14.525 -61.545 14.625 -61.445 ;
      RECT 14.525 -56.965 14.625 -56.865 ;
      RECT 14.525 -56.425 14.625 -56.325 ;
      RECT 14.525 -56.185 14.625 -56.085 ;
      RECT 14.525 -55.945 14.625 -55.845 ;
      RECT 14.525 -55.705 14.625 -55.605 ;
      RECT 14.275 -57.245 14.375 -57.145 ;
      RECT 14.275 -53.195 14.375 -53.095 ;
      RECT 14.275 -52.955 14.375 -52.855 ;
      RECT 14.275 -52.715 14.375 -52.615 ;
      RECT 14.275 -52.475 14.375 -52.375 ;
      RECT 14.015 -53.195 14.115 -53.095 ;
      RECT 14.015 -52.955 14.115 -52.855 ;
      RECT 14.015 -52.715 14.115 -52.615 ;
      RECT 14.015 -52.475 14.115 -52.375 ;
      RECT 14.015 -48.5 14.115 -48.4 ;
      RECT 14.015 -45.27 14.115 -45.17 ;
      RECT 14.015 -42.04 14.115 -41.94 ;
      RECT 14.015 -38.81 14.115 -38.71 ;
      RECT 14.015 -35.58 14.115 -35.48 ;
      RECT 14.015 -32.35 14.115 -32.25 ;
      RECT 14.015 -29.12 14.115 -29.02 ;
      RECT 14.015 -25.89 14.115 -25.79 ;
      RECT 14.015 -22.66 14.115 -22.56 ;
      RECT 14.015 -19.43 14.115 -19.33 ;
      RECT 14.015 -16.2 14.115 -16.1 ;
      RECT 14.015 -12.97 14.115 -12.87 ;
      RECT 14.015 -9.74 14.115 -9.64 ;
      RECT 14.015 -6.51 14.115 -6.41 ;
      RECT 14.015 -3.28 14.115 -3.18 ;
      RECT 14.015 -0.05 14.115 0.05 ;
      RECT 14.015 2.245 14.115 2.345 ;
      RECT 14.015 2.485 14.115 2.585 ;
      RECT 14.015 2.725 14.115 2.825 ;
      RECT 14.015 2.965 14.115 3.065 ;
      RECT 13.725 -60.485 13.825 -60.385 ;
      RECT 13.725 -60.285 13.825 -60.185 ;
      RECT 13.725 -59.015 13.825 -58.915 ;
      RECT 13.585 -53.195 13.685 -53.095 ;
      RECT 13.585 -52.955 13.685 -52.855 ;
      RECT 13.585 -52.715 13.685 -52.615 ;
      RECT 13.585 -52.475 13.685 -52.375 ;
      RECT 13.585 -48.5 13.685 -48.4 ;
      RECT 13.585 -45.27 13.685 -45.17 ;
      RECT 13.585 -42.04 13.685 -41.94 ;
      RECT 13.585 -38.81 13.685 -38.71 ;
      RECT 13.585 -35.58 13.685 -35.48 ;
      RECT 13.585 -32.35 13.685 -32.25 ;
      RECT 13.585 -29.12 13.685 -29.02 ;
      RECT 13.585 -25.89 13.685 -25.79 ;
      RECT 13.585 -22.66 13.685 -22.56 ;
      RECT 13.585 -19.43 13.685 -19.33 ;
      RECT 13.585 -16.2 13.685 -16.1 ;
      RECT 13.585 -12.97 13.685 -12.87 ;
      RECT 13.585 -9.74 13.685 -9.64 ;
      RECT 13.585 -6.51 13.685 -6.41 ;
      RECT 13.585 -3.28 13.685 -3.18 ;
      RECT 13.585 -0.05 13.685 0.05 ;
      RECT 13.585 2.245 13.685 2.345 ;
      RECT 13.585 2.485 13.685 2.585 ;
      RECT 13.585 2.725 13.685 2.825 ;
      RECT 13.585 2.965 13.685 3.065 ;
      RECT 13.325 -56.965 13.425 -56.865 ;
      RECT 13.325 -53.195 13.425 -53.095 ;
      RECT 13.325 -52.955 13.425 -52.855 ;
      RECT 13.325 -52.715 13.425 -52.615 ;
      RECT 13.325 -52.475 13.425 -52.375 ;
      RECT 13.135 -60.265 13.235 -60.165 ;
      RECT 13.135 -60.005 13.235 -59.905 ;
      RECT 13.135 -59.03 13.235 -58.93 ;
      RECT 13.135 -58.83 13.235 -58.73 ;
      RECT 13.075 -57.245 13.175 -57.145 ;
      RECT 13.075 -53.195 13.175 -53.095 ;
      RECT 13.075 -52.955 13.175 -52.855 ;
      RECT 13.075 -52.715 13.175 -52.615 ;
      RECT 13.075 -52.475 13.175 -52.375 ;
      RECT 12.835 -57.47 12.935 -57.37 ;
      RECT 12.835 -56.965 12.935 -56.865 ;
      RECT 12.815 -53.195 12.915 -53.095 ;
      RECT 12.815 -52.955 12.915 -52.855 ;
      RECT 12.815 -52.715 12.915 -52.615 ;
      RECT 12.815 -52.475 12.915 -52.375 ;
      RECT 12.815 -48.5 12.915 -48.4 ;
      RECT 12.815 -45.27 12.915 -45.17 ;
      RECT 12.815 -42.04 12.915 -41.94 ;
      RECT 12.815 -38.81 12.915 -38.71 ;
      RECT 12.815 -35.58 12.915 -35.48 ;
      RECT 12.815 -32.35 12.915 -32.25 ;
      RECT 12.815 -29.12 12.915 -29.02 ;
      RECT 12.815 -25.89 12.915 -25.79 ;
      RECT 12.815 -22.66 12.915 -22.56 ;
      RECT 12.815 -19.43 12.915 -19.33 ;
      RECT 12.815 -16.2 12.915 -16.1 ;
      RECT 12.815 -12.97 12.915 -12.87 ;
      RECT 12.815 -9.74 12.915 -9.64 ;
      RECT 12.815 -6.51 12.915 -6.41 ;
      RECT 12.815 -3.28 12.915 -3.18 ;
      RECT 12.815 -0.05 12.915 0.05 ;
      RECT 12.815 2.245 12.915 2.345 ;
      RECT 12.815 2.485 12.915 2.585 ;
      RECT 12.815 2.725 12.915 2.825 ;
      RECT 12.815 2.965 12.915 3.065 ;
      RECT 12.565 -57.875 12.665 -57.775 ;
      RECT 12.385 -53.195 12.485 -53.095 ;
      RECT 12.385 -52.955 12.485 -52.855 ;
      RECT 12.385 -52.715 12.485 -52.615 ;
      RECT 12.385 -52.475 12.485 -52.375 ;
      RECT 12.385 -48.5 12.485 -48.4 ;
      RECT 12.385 -45.27 12.485 -45.17 ;
      RECT 12.385 -42.04 12.485 -41.94 ;
      RECT 12.385 -38.81 12.485 -38.71 ;
      RECT 12.385 -35.58 12.485 -35.48 ;
      RECT 12.385 -32.35 12.485 -32.25 ;
      RECT 12.385 -29.12 12.485 -29.02 ;
      RECT 12.385 -25.89 12.485 -25.79 ;
      RECT 12.385 -22.66 12.485 -22.56 ;
      RECT 12.385 -19.43 12.485 -19.33 ;
      RECT 12.385 -16.2 12.485 -16.1 ;
      RECT 12.385 -12.97 12.485 -12.87 ;
      RECT 12.385 -9.74 12.485 -9.64 ;
      RECT 12.385 -6.51 12.485 -6.41 ;
      RECT 12.385 -3.28 12.485 -3.18 ;
      RECT 12.385 -0.05 12.485 0.05 ;
      RECT 12.385 2.245 12.485 2.345 ;
      RECT 12.385 2.485 12.485 2.585 ;
      RECT 12.385 2.725 12.485 2.825 ;
      RECT 12.385 2.965 12.485 3.065 ;
      RECT 12.24 -57.875 12.34 -57.775 ;
      RECT 12.125 -56.965 12.225 -56.865 ;
      RECT 12.125 -53.195 12.225 -53.095 ;
      RECT 12.125 -52.955 12.225 -52.855 ;
      RECT 12.125 -52.715 12.225 -52.615 ;
      RECT 12.125 -52.475 12.225 -52.375 ;
      RECT 11.875 -57.245 11.975 -57.145 ;
      RECT 11.875 -56.425 11.975 -56.325 ;
      RECT 11.875 -56.185 11.975 -56.085 ;
      RECT 11.875 -55.945 11.975 -55.845 ;
      RECT 11.875 -55.705 11.975 -55.605 ;
      RECT 11.705 -60.485 11.805 -60.385 ;
      RECT 11.705 -60.285 11.805 -60.185 ;
      RECT 11.705 -59.015 11.805 -58.915 ;
      RECT 11.615 -56.425 11.715 -56.325 ;
      RECT 11.615 -56.185 11.715 -56.085 ;
      RECT 11.615 -55.945 11.715 -55.845 ;
      RECT 11.615 -55.705 11.715 -55.605 ;
      RECT 11.615 -48.5 11.715 -48.4 ;
      RECT 11.615 -45.27 11.715 -45.17 ;
      RECT 11.615 -42.04 11.715 -41.94 ;
      RECT 11.615 -38.81 11.715 -38.71 ;
      RECT 11.615 -35.58 11.715 -35.48 ;
      RECT 11.615 -32.35 11.715 -32.25 ;
      RECT 11.615 -29.12 11.715 -29.02 ;
      RECT 11.615 -25.89 11.715 -25.79 ;
      RECT 11.615 -22.66 11.715 -22.56 ;
      RECT 11.615 -19.43 11.715 -19.33 ;
      RECT 11.615 -16.2 11.715 -16.1 ;
      RECT 11.615 -12.97 11.715 -12.87 ;
      RECT 11.615 -9.74 11.715 -9.64 ;
      RECT 11.615 -6.51 11.715 -6.41 ;
      RECT 11.615 -3.28 11.715 -3.18 ;
      RECT 11.615 -0.05 11.715 0.05 ;
      RECT 11.615 2.245 11.715 2.345 ;
      RECT 11.615 2.485 11.715 2.585 ;
      RECT 11.615 2.725 11.715 2.825 ;
      RECT 11.615 2.965 11.715 3.065 ;
      RECT 11.185 -56.425 11.285 -56.325 ;
      RECT 11.185 -56.185 11.285 -56.085 ;
      RECT 11.185 -55.945 11.285 -55.845 ;
      RECT 11.185 -55.705 11.285 -55.605 ;
      RECT 11.185 -48.5 11.285 -48.4 ;
      RECT 11.185 -45.27 11.285 -45.17 ;
      RECT 11.185 -42.04 11.285 -41.94 ;
      RECT 11.185 -38.81 11.285 -38.71 ;
      RECT 11.185 -35.58 11.285 -35.48 ;
      RECT 11.185 -32.35 11.285 -32.25 ;
      RECT 11.185 -29.12 11.285 -29.02 ;
      RECT 11.185 -25.89 11.285 -25.79 ;
      RECT 11.185 -22.66 11.285 -22.56 ;
      RECT 11.185 -19.43 11.285 -19.33 ;
      RECT 11.185 -16.2 11.285 -16.1 ;
      RECT 11.185 -12.97 11.285 -12.87 ;
      RECT 11.185 -9.74 11.285 -9.64 ;
      RECT 11.185 -6.51 11.285 -6.41 ;
      RECT 11.185 -3.28 11.285 -3.18 ;
      RECT 11.185 -0.05 11.285 0.05 ;
      RECT 11.185 2.245 11.285 2.345 ;
      RECT 11.185 2.485 11.285 2.585 ;
      RECT 11.185 2.725 11.285 2.825 ;
      RECT 11.185 2.965 11.285 3.065 ;
      RECT 11.115 -60.265 11.215 -60.165 ;
      RECT 11.115 -60.005 11.215 -59.905 ;
      RECT 11.115 -59.045 11.215 -58.945 ;
      RECT 11.115 -58.845 11.215 -58.745 ;
      RECT 10.925 -56.965 11.025 -56.865 ;
      RECT 10.925 -56.425 11.025 -56.325 ;
      RECT 10.925 -56.185 11.025 -56.085 ;
      RECT 10.925 -55.945 11.025 -55.845 ;
      RECT 10.925 -55.705 11.025 -55.605 ;
      RECT 10.675 -57.245 10.775 -57.145 ;
      RECT 10.675 -56.425 10.775 -56.325 ;
      RECT 10.675 -56.185 10.775 -56.085 ;
      RECT 10.675 -55.945 10.775 -55.845 ;
      RECT 10.675 -55.705 10.775 -55.605 ;
      RECT 10.415 -56.425 10.515 -56.325 ;
      RECT 10.415 -56.185 10.515 -56.085 ;
      RECT 10.415 -55.945 10.515 -55.845 ;
      RECT 10.415 -55.705 10.515 -55.605 ;
      RECT 10.415 -48.5 10.515 -48.4 ;
      RECT 10.415 -45.27 10.515 -45.17 ;
      RECT 10.415 -42.04 10.515 -41.94 ;
      RECT 10.415 -38.81 10.515 -38.71 ;
      RECT 10.415 -35.58 10.515 -35.48 ;
      RECT 10.415 -32.35 10.515 -32.25 ;
      RECT 10.415 -29.12 10.515 -29.02 ;
      RECT 10.415 -25.89 10.515 -25.79 ;
      RECT 10.415 -22.66 10.515 -22.56 ;
      RECT 10.415 -19.43 10.515 -19.33 ;
      RECT 10.415 -16.2 10.515 -16.1 ;
      RECT 10.415 -12.97 10.515 -12.87 ;
      RECT 10.415 -9.74 10.515 -9.64 ;
      RECT 10.415 -6.51 10.515 -6.41 ;
      RECT 10.415 -3.28 10.515 -3.18 ;
      RECT 10.415 -0.05 10.515 0.05 ;
      RECT 10.415 2.245 10.515 2.345 ;
      RECT 10.415 2.485 10.515 2.585 ;
      RECT 10.415 2.725 10.515 2.825 ;
      RECT 10.415 2.965 10.515 3.065 ;
      RECT 10.315 -61.745 10.415 -61.645 ;
      RECT 10.315 -61.545 10.415 -61.445 ;
      RECT 9.985 -56.425 10.085 -56.325 ;
      RECT 9.985 -56.185 10.085 -56.085 ;
      RECT 9.985 -55.945 10.085 -55.845 ;
      RECT 9.985 -55.705 10.085 -55.605 ;
      RECT 9.985 -48.5 10.085 -48.4 ;
      RECT 9.985 -45.27 10.085 -45.17 ;
      RECT 9.985 -42.04 10.085 -41.94 ;
      RECT 9.985 -38.81 10.085 -38.71 ;
      RECT 9.985 -35.58 10.085 -35.48 ;
      RECT 9.985 -32.35 10.085 -32.25 ;
      RECT 9.985 -29.12 10.085 -29.02 ;
      RECT 9.985 -25.89 10.085 -25.79 ;
      RECT 9.985 -22.66 10.085 -22.56 ;
      RECT 9.985 -19.43 10.085 -19.33 ;
      RECT 9.985 -16.2 10.085 -16.1 ;
      RECT 9.985 -12.97 10.085 -12.87 ;
      RECT 9.985 -9.74 10.085 -9.64 ;
      RECT 9.985 -6.51 10.085 -6.41 ;
      RECT 9.985 -3.28 10.085 -3.18 ;
      RECT 9.985 -0.05 10.085 0.05 ;
      RECT 9.985 2.245 10.085 2.345 ;
      RECT 9.985 2.485 10.085 2.585 ;
      RECT 9.985 2.725 10.085 2.825 ;
      RECT 9.985 2.965 10.085 3.065 ;
      RECT 9.965 -60.265 10.065 -60.165 ;
      RECT 9.965 -59.815 10.065 -59.715 ;
      RECT 9.965 -59.015 10.065 -58.915 ;
      RECT 9.725 -61.745 9.825 -61.645 ;
      RECT 9.725 -61.545 9.825 -61.445 ;
      RECT 9.725 -56.965 9.825 -56.865 ;
      RECT 9.725 -56.425 9.825 -56.325 ;
      RECT 9.725 -56.185 9.825 -56.085 ;
      RECT 9.725 -55.945 9.825 -55.845 ;
      RECT 9.725 -55.705 9.825 -55.605 ;
      RECT 9.475 -57.245 9.575 -57.145 ;
      RECT 9.475 -53.195 9.575 -53.095 ;
      RECT 9.475 -52.955 9.575 -52.855 ;
      RECT 9.475 -52.715 9.575 -52.615 ;
      RECT 9.475 -52.475 9.575 -52.375 ;
      RECT 9.215 -53.195 9.315 -53.095 ;
      RECT 9.215 -52.955 9.315 -52.855 ;
      RECT 9.215 -52.715 9.315 -52.615 ;
      RECT 9.215 -52.475 9.315 -52.375 ;
      RECT 9.215 -48.5 9.315 -48.4 ;
      RECT 9.215 -45.27 9.315 -45.17 ;
      RECT 9.215 -42.04 9.315 -41.94 ;
      RECT 9.215 -38.81 9.315 -38.71 ;
      RECT 9.215 -35.58 9.315 -35.48 ;
      RECT 9.215 -32.35 9.315 -32.25 ;
      RECT 9.215 -29.12 9.315 -29.02 ;
      RECT 9.215 -25.89 9.315 -25.79 ;
      RECT 9.215 -22.66 9.315 -22.56 ;
      RECT 9.215 -19.43 9.315 -19.33 ;
      RECT 9.215 -16.2 9.315 -16.1 ;
      RECT 9.215 -12.97 9.315 -12.87 ;
      RECT 9.215 -9.74 9.315 -9.64 ;
      RECT 9.215 -6.51 9.315 -6.41 ;
      RECT 9.215 -3.28 9.315 -3.18 ;
      RECT 9.215 -0.05 9.315 0.05 ;
      RECT 9.215 2.245 9.315 2.345 ;
      RECT 9.215 2.485 9.315 2.585 ;
      RECT 9.215 2.725 9.315 2.825 ;
      RECT 9.215 2.965 9.315 3.065 ;
      RECT 8.925 -60.485 9.025 -60.385 ;
      RECT 8.925 -60.285 9.025 -60.185 ;
      RECT 8.925 -59.015 9.025 -58.915 ;
      RECT 8.785 -53.195 8.885 -53.095 ;
      RECT 8.785 -52.955 8.885 -52.855 ;
      RECT 8.785 -52.715 8.885 -52.615 ;
      RECT 8.785 -52.475 8.885 -52.375 ;
      RECT 8.785 -48.5 8.885 -48.4 ;
      RECT 8.785 -45.27 8.885 -45.17 ;
      RECT 8.785 -42.04 8.885 -41.94 ;
      RECT 8.785 -38.81 8.885 -38.71 ;
      RECT 8.785 -35.58 8.885 -35.48 ;
      RECT 8.785 -32.35 8.885 -32.25 ;
      RECT 8.785 -29.12 8.885 -29.02 ;
      RECT 8.785 -25.89 8.885 -25.79 ;
      RECT 8.785 -22.66 8.885 -22.56 ;
      RECT 8.785 -19.43 8.885 -19.33 ;
      RECT 8.785 -16.2 8.885 -16.1 ;
      RECT 8.785 -12.97 8.885 -12.87 ;
      RECT 8.785 -9.74 8.885 -9.64 ;
      RECT 8.785 -6.51 8.885 -6.41 ;
      RECT 8.785 -3.28 8.885 -3.18 ;
      RECT 8.785 -0.05 8.885 0.05 ;
      RECT 8.785 2.245 8.885 2.345 ;
      RECT 8.785 2.485 8.885 2.585 ;
      RECT 8.785 2.725 8.885 2.825 ;
      RECT 8.785 2.965 8.885 3.065 ;
      RECT 8.525 -56.965 8.625 -56.865 ;
      RECT 8.525 -53.195 8.625 -53.095 ;
      RECT 8.525 -52.955 8.625 -52.855 ;
      RECT 8.525 -52.715 8.625 -52.615 ;
      RECT 8.525 -52.475 8.625 -52.375 ;
      RECT 8.335 -60.265 8.435 -60.165 ;
      RECT 8.335 -60.005 8.435 -59.905 ;
      RECT 8.335 -59.03 8.435 -58.93 ;
      RECT 8.335 -58.83 8.435 -58.73 ;
      RECT 8.275 -57.245 8.375 -57.145 ;
      RECT 8.275 -53.195 8.375 -53.095 ;
      RECT 8.275 -52.955 8.375 -52.855 ;
      RECT 8.275 -52.715 8.375 -52.615 ;
      RECT 8.275 -52.475 8.375 -52.375 ;
      RECT 8.035 -57.47 8.135 -57.37 ;
      RECT 8.035 -56.965 8.135 -56.865 ;
      RECT 8.015 -53.195 8.115 -53.095 ;
      RECT 8.015 -52.955 8.115 -52.855 ;
      RECT 8.015 -52.715 8.115 -52.615 ;
      RECT 8.015 -52.475 8.115 -52.375 ;
      RECT 8.015 -48.5 8.115 -48.4 ;
      RECT 8.015 -45.27 8.115 -45.17 ;
      RECT 8.015 -42.04 8.115 -41.94 ;
      RECT 8.015 -38.81 8.115 -38.71 ;
      RECT 8.015 -35.58 8.115 -35.48 ;
      RECT 8.015 -32.35 8.115 -32.25 ;
      RECT 8.015 -29.12 8.115 -29.02 ;
      RECT 8.015 -25.89 8.115 -25.79 ;
      RECT 8.015 -22.66 8.115 -22.56 ;
      RECT 8.015 -19.43 8.115 -19.33 ;
      RECT 8.015 -16.2 8.115 -16.1 ;
      RECT 8.015 -12.97 8.115 -12.87 ;
      RECT 8.015 -9.74 8.115 -9.64 ;
      RECT 8.015 -6.51 8.115 -6.41 ;
      RECT 8.015 -3.28 8.115 -3.18 ;
      RECT 8.015 -0.05 8.115 0.05 ;
      RECT 8.015 2.245 8.115 2.345 ;
      RECT 8.015 2.485 8.115 2.585 ;
      RECT 8.015 2.725 8.115 2.825 ;
      RECT 8.015 2.965 8.115 3.065 ;
      RECT 7.765 -57.875 7.865 -57.775 ;
      RECT 7.585 -53.195 7.685 -53.095 ;
      RECT 7.585 -52.955 7.685 -52.855 ;
      RECT 7.585 -52.715 7.685 -52.615 ;
      RECT 7.585 -52.475 7.685 -52.375 ;
      RECT 7.585 -48.5 7.685 -48.4 ;
      RECT 7.585 -45.27 7.685 -45.17 ;
      RECT 7.585 -42.04 7.685 -41.94 ;
      RECT 7.585 -38.81 7.685 -38.71 ;
      RECT 7.585 -35.58 7.685 -35.48 ;
      RECT 7.585 -32.35 7.685 -32.25 ;
      RECT 7.585 -29.12 7.685 -29.02 ;
      RECT 7.585 -25.89 7.685 -25.79 ;
      RECT 7.585 -22.66 7.685 -22.56 ;
      RECT 7.585 -19.43 7.685 -19.33 ;
      RECT 7.585 -16.2 7.685 -16.1 ;
      RECT 7.585 -12.97 7.685 -12.87 ;
      RECT 7.585 -9.74 7.685 -9.64 ;
      RECT 7.585 -6.51 7.685 -6.41 ;
      RECT 7.585 -3.28 7.685 -3.18 ;
      RECT 7.585 -0.05 7.685 0.05 ;
      RECT 7.585 2.245 7.685 2.345 ;
      RECT 7.585 2.485 7.685 2.585 ;
      RECT 7.585 2.725 7.685 2.825 ;
      RECT 7.585 2.965 7.685 3.065 ;
      RECT 7.44 -57.875 7.54 -57.775 ;
      RECT 7.325 -56.965 7.425 -56.865 ;
      RECT 7.325 -53.195 7.425 -53.095 ;
      RECT 7.325 -52.955 7.425 -52.855 ;
      RECT 7.325 -52.715 7.425 -52.615 ;
      RECT 7.325 -52.475 7.425 -52.375 ;
      RECT 7.075 -57.245 7.175 -57.145 ;
      RECT 7.075 -56.425 7.175 -56.325 ;
      RECT 7.075 -56.185 7.175 -56.085 ;
      RECT 7.075 -55.945 7.175 -55.845 ;
      RECT 7.075 -55.705 7.175 -55.605 ;
      RECT 6.905 -60.485 7.005 -60.385 ;
      RECT 6.905 -60.285 7.005 -60.185 ;
      RECT 6.905 -59.015 7.005 -58.915 ;
      RECT 6.815 -56.425 6.915 -56.325 ;
      RECT 6.815 -56.185 6.915 -56.085 ;
      RECT 6.815 -55.945 6.915 -55.845 ;
      RECT 6.815 -55.705 6.915 -55.605 ;
      RECT 6.815 -48.5 6.915 -48.4 ;
      RECT 6.815 -45.27 6.915 -45.17 ;
      RECT 6.815 -42.04 6.915 -41.94 ;
      RECT 6.815 -38.81 6.915 -38.71 ;
      RECT 6.815 -35.58 6.915 -35.48 ;
      RECT 6.815 -32.35 6.915 -32.25 ;
      RECT 6.815 -29.12 6.915 -29.02 ;
      RECT 6.815 -25.89 6.915 -25.79 ;
      RECT 6.815 -22.66 6.915 -22.56 ;
      RECT 6.815 -19.43 6.915 -19.33 ;
      RECT 6.815 -16.2 6.915 -16.1 ;
      RECT 6.815 -12.97 6.915 -12.87 ;
      RECT 6.815 -9.74 6.915 -9.64 ;
      RECT 6.815 -6.51 6.915 -6.41 ;
      RECT 6.815 -3.28 6.915 -3.18 ;
      RECT 6.815 -0.05 6.915 0.05 ;
      RECT 6.815 2.245 6.915 2.345 ;
      RECT 6.815 2.485 6.915 2.585 ;
      RECT 6.815 2.725 6.915 2.825 ;
      RECT 6.815 2.965 6.915 3.065 ;
      RECT 6.385 -56.425 6.485 -56.325 ;
      RECT 6.385 -56.185 6.485 -56.085 ;
      RECT 6.385 -55.945 6.485 -55.845 ;
      RECT 6.385 -55.705 6.485 -55.605 ;
      RECT 6.385 -48.5 6.485 -48.4 ;
      RECT 6.385 -45.27 6.485 -45.17 ;
      RECT 6.385 -42.04 6.485 -41.94 ;
      RECT 6.385 -38.81 6.485 -38.71 ;
      RECT 6.385 -35.58 6.485 -35.48 ;
      RECT 6.385 -32.35 6.485 -32.25 ;
      RECT 6.385 -29.12 6.485 -29.02 ;
      RECT 6.385 -25.89 6.485 -25.79 ;
      RECT 6.385 -22.66 6.485 -22.56 ;
      RECT 6.385 -19.43 6.485 -19.33 ;
      RECT 6.385 -16.2 6.485 -16.1 ;
      RECT 6.385 -12.97 6.485 -12.87 ;
      RECT 6.385 -9.74 6.485 -9.64 ;
      RECT 6.385 -6.51 6.485 -6.41 ;
      RECT 6.385 -3.28 6.485 -3.18 ;
      RECT 6.385 -0.05 6.485 0.05 ;
      RECT 6.385 2.245 6.485 2.345 ;
      RECT 6.385 2.485 6.485 2.585 ;
      RECT 6.385 2.725 6.485 2.825 ;
      RECT 6.385 2.965 6.485 3.065 ;
      RECT 6.315 -60.265 6.415 -60.165 ;
      RECT 6.315 -60.005 6.415 -59.905 ;
      RECT 6.315 -59.045 6.415 -58.945 ;
      RECT 6.315 -58.845 6.415 -58.745 ;
      RECT 6.125 -56.965 6.225 -56.865 ;
      RECT 6.125 -56.425 6.225 -56.325 ;
      RECT 6.125 -56.185 6.225 -56.085 ;
      RECT 6.125 -55.945 6.225 -55.845 ;
      RECT 6.125 -55.705 6.225 -55.605 ;
      RECT 5.875 -57.245 5.975 -57.145 ;
      RECT 5.875 -56.425 5.975 -56.325 ;
      RECT 5.875 -56.185 5.975 -56.085 ;
      RECT 5.875 -55.945 5.975 -55.845 ;
      RECT 5.875 -55.705 5.975 -55.605 ;
      RECT 5.615 -56.425 5.715 -56.325 ;
      RECT 5.615 -56.185 5.715 -56.085 ;
      RECT 5.615 -55.945 5.715 -55.845 ;
      RECT 5.615 -55.705 5.715 -55.605 ;
      RECT 5.615 -48.5 5.715 -48.4 ;
      RECT 5.615 -45.27 5.715 -45.17 ;
      RECT 5.615 -42.04 5.715 -41.94 ;
      RECT 5.615 -38.81 5.715 -38.71 ;
      RECT 5.615 -35.58 5.715 -35.48 ;
      RECT 5.615 -32.35 5.715 -32.25 ;
      RECT 5.615 -29.12 5.715 -29.02 ;
      RECT 5.615 -25.89 5.715 -25.79 ;
      RECT 5.615 -22.66 5.715 -22.56 ;
      RECT 5.615 -19.43 5.715 -19.33 ;
      RECT 5.615 -16.2 5.715 -16.1 ;
      RECT 5.615 -12.97 5.715 -12.87 ;
      RECT 5.615 -9.74 5.715 -9.64 ;
      RECT 5.615 -6.51 5.715 -6.41 ;
      RECT 5.615 -3.28 5.715 -3.18 ;
      RECT 5.615 -0.05 5.715 0.05 ;
      RECT 5.615 2.245 5.715 2.345 ;
      RECT 5.615 2.485 5.715 2.585 ;
      RECT 5.615 2.725 5.715 2.825 ;
      RECT 5.615 2.965 5.715 3.065 ;
      RECT 5.515 -61.745 5.615 -61.645 ;
      RECT 5.515 -61.545 5.615 -61.445 ;
      RECT 5.185 -56.425 5.285 -56.325 ;
      RECT 5.185 -56.185 5.285 -56.085 ;
      RECT 5.185 -55.945 5.285 -55.845 ;
      RECT 5.185 -55.705 5.285 -55.605 ;
      RECT 5.185 -48.5 5.285 -48.4 ;
      RECT 5.185 -45.27 5.285 -45.17 ;
      RECT 5.185 -42.04 5.285 -41.94 ;
      RECT 5.185 -38.81 5.285 -38.71 ;
      RECT 5.185 -35.58 5.285 -35.48 ;
      RECT 5.185 -32.35 5.285 -32.25 ;
      RECT 5.185 -29.12 5.285 -29.02 ;
      RECT 5.185 -25.89 5.285 -25.79 ;
      RECT 5.185 -22.66 5.285 -22.56 ;
      RECT 5.185 -19.43 5.285 -19.33 ;
      RECT 5.185 -16.2 5.285 -16.1 ;
      RECT 5.185 -12.97 5.285 -12.87 ;
      RECT 5.185 -9.74 5.285 -9.64 ;
      RECT 5.185 -6.51 5.285 -6.41 ;
      RECT 5.185 -3.28 5.285 -3.18 ;
      RECT 5.185 -0.05 5.285 0.05 ;
      RECT 5.185 2.245 5.285 2.345 ;
      RECT 5.185 2.485 5.285 2.585 ;
      RECT 5.185 2.725 5.285 2.825 ;
      RECT 5.185 2.965 5.285 3.065 ;
      RECT 5.165 -60.265 5.265 -60.165 ;
      RECT 5.165 -59.815 5.265 -59.715 ;
      RECT 5.165 -59.015 5.265 -58.915 ;
      RECT 4.925 -61.745 5.025 -61.645 ;
      RECT 4.925 -61.545 5.025 -61.445 ;
      RECT 4.925 -56.965 5.025 -56.865 ;
      RECT 4.925 -56.425 5.025 -56.325 ;
      RECT 4.925 -56.185 5.025 -56.085 ;
      RECT 4.925 -55.945 5.025 -55.845 ;
      RECT 4.925 -55.705 5.025 -55.605 ;
      RECT 4.675 -57.245 4.775 -57.145 ;
      RECT 4.675 -53.195 4.775 -53.095 ;
      RECT 4.675 -52.955 4.775 -52.855 ;
      RECT 4.675 -52.715 4.775 -52.615 ;
      RECT 4.675 -52.475 4.775 -52.375 ;
      RECT 4.415 -53.195 4.515 -53.095 ;
      RECT 4.415 -52.955 4.515 -52.855 ;
      RECT 4.415 -52.715 4.515 -52.615 ;
      RECT 4.415 -52.475 4.515 -52.375 ;
      RECT 4.415 -48.5 4.515 -48.4 ;
      RECT 4.415 -45.27 4.515 -45.17 ;
      RECT 4.415 -42.04 4.515 -41.94 ;
      RECT 4.415 -38.81 4.515 -38.71 ;
      RECT 4.415 -35.58 4.515 -35.48 ;
      RECT 4.415 -32.35 4.515 -32.25 ;
      RECT 4.415 -29.12 4.515 -29.02 ;
      RECT 4.415 -25.89 4.515 -25.79 ;
      RECT 4.415 -22.66 4.515 -22.56 ;
      RECT 4.415 -19.43 4.515 -19.33 ;
      RECT 4.415 -16.2 4.515 -16.1 ;
      RECT 4.415 -12.97 4.515 -12.87 ;
      RECT 4.415 -9.74 4.515 -9.64 ;
      RECT 4.415 -6.51 4.515 -6.41 ;
      RECT 4.415 -3.28 4.515 -3.18 ;
      RECT 4.415 -0.05 4.515 0.05 ;
      RECT 4.415 2.245 4.515 2.345 ;
      RECT 4.415 2.485 4.515 2.585 ;
      RECT 4.415 2.725 4.515 2.825 ;
      RECT 4.415 2.965 4.515 3.065 ;
      RECT 4.125 -60.485 4.225 -60.385 ;
      RECT 4.125 -60.285 4.225 -60.185 ;
      RECT 4.125 -59.015 4.225 -58.915 ;
      RECT 3.985 -53.195 4.085 -53.095 ;
      RECT 3.985 -52.955 4.085 -52.855 ;
      RECT 3.985 -52.715 4.085 -52.615 ;
      RECT 3.985 -52.475 4.085 -52.375 ;
      RECT 3.985 -48.5 4.085 -48.4 ;
      RECT 3.985 -45.27 4.085 -45.17 ;
      RECT 3.985 -42.04 4.085 -41.94 ;
      RECT 3.985 -38.81 4.085 -38.71 ;
      RECT 3.985 -35.58 4.085 -35.48 ;
      RECT 3.985 -32.35 4.085 -32.25 ;
      RECT 3.985 -29.12 4.085 -29.02 ;
      RECT 3.985 -25.89 4.085 -25.79 ;
      RECT 3.985 -22.66 4.085 -22.56 ;
      RECT 3.985 -19.43 4.085 -19.33 ;
      RECT 3.985 -16.2 4.085 -16.1 ;
      RECT 3.985 -12.97 4.085 -12.87 ;
      RECT 3.985 -9.74 4.085 -9.64 ;
      RECT 3.985 -6.51 4.085 -6.41 ;
      RECT 3.985 -3.28 4.085 -3.18 ;
      RECT 3.985 -0.05 4.085 0.05 ;
      RECT 3.985 2.245 4.085 2.345 ;
      RECT 3.985 2.485 4.085 2.585 ;
      RECT 3.985 2.725 4.085 2.825 ;
      RECT 3.985 2.965 4.085 3.065 ;
      RECT 3.725 -56.965 3.825 -56.865 ;
      RECT 3.725 -53.195 3.825 -53.095 ;
      RECT 3.725 -52.955 3.825 -52.855 ;
      RECT 3.725 -52.715 3.825 -52.615 ;
      RECT 3.725 -52.475 3.825 -52.375 ;
      RECT 3.535 -60.265 3.635 -60.165 ;
      RECT 3.535 -60.005 3.635 -59.905 ;
      RECT 3.535 -59.03 3.635 -58.93 ;
      RECT 3.535 -58.83 3.635 -58.73 ;
      RECT 3.475 -57.245 3.575 -57.145 ;
      RECT 3.475 -53.195 3.575 -53.095 ;
      RECT 3.475 -52.955 3.575 -52.855 ;
      RECT 3.475 -52.715 3.575 -52.615 ;
      RECT 3.475 -52.475 3.575 -52.375 ;
      RECT 3.235 -57.47 3.335 -57.37 ;
      RECT 3.235 -56.965 3.335 -56.865 ;
      RECT 3.215 -53.195 3.315 -53.095 ;
      RECT 3.215 -52.955 3.315 -52.855 ;
      RECT 3.215 -52.715 3.315 -52.615 ;
      RECT 3.215 -52.475 3.315 -52.375 ;
      RECT 3.215 -48.5 3.315 -48.4 ;
      RECT 3.215 -45.27 3.315 -45.17 ;
      RECT 3.215 -42.04 3.315 -41.94 ;
      RECT 3.215 -38.81 3.315 -38.71 ;
      RECT 3.215 -35.58 3.315 -35.48 ;
      RECT 3.215 -32.35 3.315 -32.25 ;
      RECT 3.215 -29.12 3.315 -29.02 ;
      RECT 3.215 -25.89 3.315 -25.79 ;
      RECT 3.215 -22.66 3.315 -22.56 ;
      RECT 3.215 -19.43 3.315 -19.33 ;
      RECT 3.215 -16.2 3.315 -16.1 ;
      RECT 3.215 -12.97 3.315 -12.87 ;
      RECT 3.215 -9.74 3.315 -9.64 ;
      RECT 3.215 -6.51 3.315 -6.41 ;
      RECT 3.215 -3.28 3.315 -3.18 ;
      RECT 3.215 -0.05 3.315 0.05 ;
      RECT 3.215 2.245 3.315 2.345 ;
      RECT 3.215 2.485 3.315 2.585 ;
      RECT 3.215 2.725 3.315 2.825 ;
      RECT 3.215 2.965 3.315 3.065 ;
      RECT 2.965 -57.875 3.065 -57.775 ;
      RECT 2.785 -53.195 2.885 -53.095 ;
      RECT 2.785 -52.955 2.885 -52.855 ;
      RECT 2.785 -52.715 2.885 -52.615 ;
      RECT 2.785 -52.475 2.885 -52.375 ;
      RECT 2.785 -48.5 2.885 -48.4 ;
      RECT 2.785 -45.27 2.885 -45.17 ;
      RECT 2.785 -42.04 2.885 -41.94 ;
      RECT 2.785 -38.81 2.885 -38.71 ;
      RECT 2.785 -35.58 2.885 -35.48 ;
      RECT 2.785 -32.35 2.885 -32.25 ;
      RECT 2.785 -29.12 2.885 -29.02 ;
      RECT 2.785 -25.89 2.885 -25.79 ;
      RECT 2.785 -22.66 2.885 -22.56 ;
      RECT 2.785 -19.43 2.885 -19.33 ;
      RECT 2.785 -16.2 2.885 -16.1 ;
      RECT 2.785 -12.97 2.885 -12.87 ;
      RECT 2.785 -9.74 2.885 -9.64 ;
      RECT 2.785 -6.51 2.885 -6.41 ;
      RECT 2.785 -3.28 2.885 -3.18 ;
      RECT 2.785 -0.05 2.885 0.05 ;
      RECT 2.785 2.245 2.885 2.345 ;
      RECT 2.785 2.485 2.885 2.585 ;
      RECT 2.785 2.725 2.885 2.825 ;
      RECT 2.785 2.965 2.885 3.065 ;
      RECT 2.64 -57.875 2.74 -57.775 ;
      RECT 2.525 -56.965 2.625 -56.865 ;
      RECT 2.525 -53.195 2.625 -53.095 ;
      RECT 2.525 -52.955 2.625 -52.855 ;
      RECT 2.525 -52.715 2.625 -52.615 ;
      RECT 2.525 -52.475 2.625 -52.375 ;
      RECT 2.275 -57.245 2.375 -57.145 ;
      RECT 2.275 -56.425 2.375 -56.325 ;
      RECT 2.275 -56.185 2.375 -56.085 ;
      RECT 2.275 -55.945 2.375 -55.845 ;
      RECT 2.275 -55.705 2.375 -55.605 ;
      RECT 2.105 -60.485 2.205 -60.385 ;
      RECT 2.105 -60.285 2.205 -60.185 ;
      RECT 2.105 -59.015 2.205 -58.915 ;
      RECT 2.015 -56.425 2.115 -56.325 ;
      RECT 2.015 -56.185 2.115 -56.085 ;
      RECT 2.015 -55.945 2.115 -55.845 ;
      RECT 2.015 -55.705 2.115 -55.605 ;
      RECT 2.015 -48.5 2.115 -48.4 ;
      RECT 2.015 -45.27 2.115 -45.17 ;
      RECT 2.015 -42.04 2.115 -41.94 ;
      RECT 2.015 -38.81 2.115 -38.71 ;
      RECT 2.015 -35.58 2.115 -35.48 ;
      RECT 2.015 -32.35 2.115 -32.25 ;
      RECT 2.015 -29.12 2.115 -29.02 ;
      RECT 2.015 -25.89 2.115 -25.79 ;
      RECT 2.015 -22.66 2.115 -22.56 ;
      RECT 2.015 -19.43 2.115 -19.33 ;
      RECT 2.015 -16.2 2.115 -16.1 ;
      RECT 2.015 -12.97 2.115 -12.87 ;
      RECT 2.015 -9.74 2.115 -9.64 ;
      RECT 2.015 -6.51 2.115 -6.41 ;
      RECT 2.015 -3.28 2.115 -3.18 ;
      RECT 2.015 -0.05 2.115 0.05 ;
      RECT 2.015 2.245 2.115 2.345 ;
      RECT 2.015 2.485 2.115 2.585 ;
      RECT 2.015 2.725 2.115 2.825 ;
      RECT 2.015 2.965 2.115 3.065 ;
      RECT 1.585 -56.425 1.685 -56.325 ;
      RECT 1.585 -56.185 1.685 -56.085 ;
      RECT 1.585 -55.945 1.685 -55.845 ;
      RECT 1.585 -55.705 1.685 -55.605 ;
      RECT 1.585 -48.5 1.685 -48.4 ;
      RECT 1.585 -45.27 1.685 -45.17 ;
      RECT 1.585 -42.04 1.685 -41.94 ;
      RECT 1.585 -38.81 1.685 -38.71 ;
      RECT 1.585 -35.58 1.685 -35.48 ;
      RECT 1.585 -32.35 1.685 -32.25 ;
      RECT 1.585 -29.12 1.685 -29.02 ;
      RECT 1.585 -25.89 1.685 -25.79 ;
      RECT 1.585 -22.66 1.685 -22.56 ;
      RECT 1.585 -19.43 1.685 -19.33 ;
      RECT 1.585 -16.2 1.685 -16.1 ;
      RECT 1.585 -12.97 1.685 -12.87 ;
      RECT 1.585 -9.74 1.685 -9.64 ;
      RECT 1.585 -6.51 1.685 -6.41 ;
      RECT 1.585 -3.28 1.685 -3.18 ;
      RECT 1.585 -0.05 1.685 0.05 ;
      RECT 1.585 2.245 1.685 2.345 ;
      RECT 1.585 2.485 1.685 2.585 ;
      RECT 1.585 2.725 1.685 2.825 ;
      RECT 1.585 2.965 1.685 3.065 ;
      RECT 1.515 -60.265 1.615 -60.165 ;
      RECT 1.515 -60.005 1.615 -59.905 ;
      RECT 1.515 -59.045 1.615 -58.945 ;
      RECT 1.515 -58.845 1.615 -58.745 ;
      RECT 1.325 -56.965 1.425 -56.865 ;
      RECT 1.325 -56.425 1.425 -56.325 ;
      RECT 1.325 -56.185 1.425 -56.085 ;
      RECT 1.325 -55.945 1.425 -55.845 ;
      RECT 1.325 -55.705 1.425 -55.605 ;
      RECT 1.075 -57.245 1.175 -57.145 ;
      RECT 1.075 -56.425 1.175 -56.325 ;
      RECT 1.075 -56.185 1.175 -56.085 ;
      RECT 1.075 -55.945 1.175 -55.845 ;
      RECT 1.075 -55.705 1.175 -55.605 ;
      RECT 0.815 -56.425 0.915 -56.325 ;
      RECT 0.815 -56.185 0.915 -56.085 ;
      RECT 0.815 -55.945 0.915 -55.845 ;
      RECT 0.815 -55.705 0.915 -55.605 ;
      RECT 0.815 -48.5 0.915 -48.4 ;
      RECT 0.815 -45.27 0.915 -45.17 ;
      RECT 0.815 -42.04 0.915 -41.94 ;
      RECT 0.815 -38.81 0.915 -38.71 ;
      RECT 0.815 -35.58 0.915 -35.48 ;
      RECT 0.815 -32.35 0.915 -32.25 ;
      RECT 0.815 -29.12 0.915 -29.02 ;
      RECT 0.815 -25.89 0.915 -25.79 ;
      RECT 0.815 -22.66 0.915 -22.56 ;
      RECT 0.815 -19.43 0.915 -19.33 ;
      RECT 0.815 -16.2 0.915 -16.1 ;
      RECT 0.815 -12.97 0.915 -12.87 ;
      RECT 0.815 -9.74 0.915 -9.64 ;
      RECT 0.815 -6.51 0.915 -6.41 ;
      RECT 0.815 -3.28 0.915 -3.18 ;
      RECT 0.815 -0.05 0.915 0.05 ;
      RECT 0.815 2.245 0.915 2.345 ;
      RECT 0.815 2.485 0.915 2.585 ;
      RECT 0.815 2.725 0.915 2.825 ;
      RECT 0.815 2.965 0.915 3.065 ;
      RECT 0.715 -61.745 0.815 -61.645 ;
      RECT 0.715 -61.545 0.815 -61.445 ;
      RECT 0.385 -56.425 0.485 -56.325 ;
      RECT 0.385 -56.185 0.485 -56.085 ;
      RECT 0.385 -55.945 0.485 -55.845 ;
      RECT 0.385 -55.705 0.485 -55.605 ;
      RECT 0.385 -48.5 0.485 -48.4 ;
      RECT 0.385 -45.27 0.485 -45.17 ;
      RECT 0.385 -42.04 0.485 -41.94 ;
      RECT 0.385 -38.81 0.485 -38.71 ;
      RECT 0.385 -35.58 0.485 -35.48 ;
      RECT 0.385 -32.35 0.485 -32.25 ;
      RECT 0.385 -29.12 0.485 -29.02 ;
      RECT 0.385 -25.89 0.485 -25.79 ;
      RECT 0.385 -22.66 0.485 -22.56 ;
      RECT 0.385 -19.43 0.485 -19.33 ;
      RECT 0.385 -16.2 0.485 -16.1 ;
      RECT 0.385 -12.97 0.485 -12.87 ;
      RECT 0.385 -9.74 0.485 -9.64 ;
      RECT 0.385 -6.51 0.485 -6.41 ;
      RECT 0.385 -3.28 0.485 -3.18 ;
      RECT 0.385 -0.05 0.485 0.05 ;
      RECT 0.385 2.245 0.485 2.345 ;
      RECT 0.385 2.485 0.485 2.585 ;
      RECT 0.385 2.725 0.485 2.825 ;
      RECT 0.385 2.965 0.485 3.065 ;
      RECT 0.365 -60.265 0.465 -60.165 ;
      RECT 0.365 -59.815 0.465 -59.715 ;
      RECT 0.365 -59.015 0.465 -58.915 ;
      RECT 0.125 -61.745 0.225 -61.645 ;
      RECT 0.125 -61.545 0.225 -61.445 ;
      RECT 0.125 -56.965 0.225 -56.865 ;
      RECT 0.125 -56.425 0.225 -56.325 ;
      RECT 0.125 -56.185 0.225 -56.085 ;
      RECT 0.125 -55.945 0.225 -55.845 ;
      RECT 0.125 -55.705 0.225 -55.605 ;
      RECT -0.385 1.935 -0.285 2.035 ;
      RECT -0.385 4.135 -0.285 4.235 ;
      RECT -0.765 -55.905 -0.665 -55.805 ;
      RECT -0.765 -55.22 -0.665 -55.12 ;
      RECT -0.765 -51.145 -0.665 -51.045 ;
      RECT -0.765 -50.905 -0.665 -50.805 ;
      RECT -0.765 -49.325 -0.665 -49.225 ;
      RECT -0.765 -49.085 -0.665 -48.985 ;
      RECT -0.765 -45.01 -0.665 -44.91 ;
      RECT -0.765 -44.325 -0.665 -44.225 ;
      RECT -0.765 -42.985 -0.665 -42.885 ;
      RECT -0.765 -42.3 -0.665 -42.2 ;
      RECT -0.765 -38.225 -0.665 -38.125 ;
      RECT -0.765 -37.985 -0.665 -37.885 ;
      RECT -0.765 -36.405 -0.665 -36.305 ;
      RECT -0.765 -36.165 -0.665 -36.065 ;
      RECT -0.765 -32.09 -0.665 -31.99 ;
      RECT -0.765 -31.405 -0.665 -31.305 ;
      RECT -0.765 -30.065 -0.665 -29.965 ;
      RECT -0.765 -29.38 -0.665 -29.28 ;
      RECT -0.765 -25.305 -0.665 -25.205 ;
      RECT -0.765 -25.065 -0.665 -24.965 ;
      RECT -0.765 -23.485 -0.665 -23.385 ;
      RECT -0.765 -23.245 -0.665 -23.145 ;
      RECT -0.765 -19.17 -0.665 -19.07 ;
      RECT -0.765 -18.485 -0.665 -18.385 ;
      RECT -0.765 -17.145 -0.665 -17.045 ;
      RECT -0.765 -16.46 -0.665 -16.36 ;
      RECT -0.765 -12.385 -0.665 -12.285 ;
      RECT -0.765 -12.145 -0.665 -12.045 ;
      RECT -0.765 -10.565 -0.665 -10.465 ;
      RECT -0.765 -10.325 -0.665 -10.225 ;
      RECT -0.765 -6.25 -0.665 -6.15 ;
      RECT -0.765 -5.565 -0.665 -5.465 ;
      RECT -0.765 -4.225 -0.665 -4.125 ;
      RECT -0.765 -3.54 -0.665 -3.44 ;
      RECT -0.765 0.535 -0.665 0.635 ;
      RECT -0.765 0.775 -0.665 0.875 ;
      RECT -1.285 -55.905 -1.185 -55.805 ;
      RECT -1.285 -55.665 -1.185 -55.565 ;
      RECT -1.285 -51.73 -1.185 -51.63 ;
      RECT -1.285 -51.145 -1.185 -51.045 ;
      RECT -1.285 -50.905 -1.185 -50.805 ;
      RECT -1.285 -49.325 -1.185 -49.225 ;
      RECT -1.285 -49.085 -1.185 -48.985 ;
      RECT -1.285 -48.5 -1.185 -48.4 ;
      RECT -1.285 -44.565 -1.185 -44.465 ;
      RECT -1.285 -44.325 -1.185 -44.225 ;
      RECT -1.285 -42.985 -1.185 -42.885 ;
      RECT -1.285 -42.745 -1.185 -42.645 ;
      RECT -1.285 -38.81 -1.185 -38.71 ;
      RECT -1.285 -38.225 -1.185 -38.125 ;
      RECT -1.285 -37.985 -1.185 -37.885 ;
      RECT -1.285 -36.405 -1.185 -36.305 ;
      RECT -1.285 -36.165 -1.185 -36.065 ;
      RECT -1.285 -35.58 -1.185 -35.48 ;
      RECT -1.285 -31.645 -1.185 -31.545 ;
      RECT -1.285 -31.405 -1.185 -31.305 ;
      RECT -1.285 -30.065 -1.185 -29.965 ;
      RECT -1.285 -29.825 -1.185 -29.725 ;
      RECT -1.285 -25.89 -1.185 -25.79 ;
      RECT -1.285 -25.305 -1.185 -25.205 ;
      RECT -1.285 -25.065 -1.185 -24.965 ;
      RECT -1.285 -23.485 -1.185 -23.385 ;
      RECT -1.285 -23.245 -1.185 -23.145 ;
      RECT -1.285 -22.66 -1.185 -22.56 ;
      RECT -1.285 -18.725 -1.185 -18.625 ;
      RECT -1.285 -18.485 -1.185 -18.385 ;
      RECT -1.285 -17.145 -1.185 -17.045 ;
      RECT -1.285 -16.905 -1.185 -16.805 ;
      RECT -1.285 -12.97 -1.185 -12.87 ;
      RECT -1.285 -12.385 -1.185 -12.285 ;
      RECT -1.285 -12.145 -1.185 -12.045 ;
      RECT -1.285 -10.565 -1.185 -10.465 ;
      RECT -1.285 -10.325 -1.185 -10.225 ;
      RECT -1.285 -9.74 -1.185 -9.64 ;
      RECT -1.285 -5.805 -1.185 -5.705 ;
      RECT -1.285 -5.565 -1.185 -5.465 ;
      RECT -1.285 -4.225 -1.185 -4.125 ;
      RECT -1.285 -3.985 -1.185 -3.885 ;
      RECT -1.285 -0.05 -1.185 0.05 ;
      RECT -1.285 0.535 -1.185 0.635 ;
      RECT -1.285 0.775 -1.185 0.875 ;
      RECT -1.805 -51.73 -1.705 -51.63 ;
      RECT -1.805 -51.145 -1.705 -51.045 ;
      RECT -1.805 -50.905 -1.705 -50.805 ;
      RECT -1.805 -49.325 -1.705 -49.225 ;
      RECT -1.805 -49.085 -1.705 -48.985 ;
      RECT -1.805 -48.5 -1.705 -48.4 ;
      RECT -1.805 -38.81 -1.705 -38.71 ;
      RECT -1.805 -38.225 -1.705 -38.125 ;
      RECT -1.805 -37.985 -1.705 -37.885 ;
      RECT -1.805 -36.405 -1.705 -36.305 ;
      RECT -1.805 -36.165 -1.705 -36.065 ;
      RECT -1.805 -35.58 -1.705 -35.48 ;
      RECT -1.805 -25.89 -1.705 -25.79 ;
      RECT -1.805 -25.305 -1.705 -25.205 ;
      RECT -1.805 -25.065 -1.705 -24.965 ;
      RECT -1.805 -23.485 -1.705 -23.385 ;
      RECT -1.805 -23.245 -1.705 -23.145 ;
      RECT -1.805 -22.66 -1.705 -22.56 ;
      RECT -1.805 -12.97 -1.705 -12.87 ;
      RECT -1.805 -12.385 -1.705 -12.285 ;
      RECT -1.805 -12.145 -1.705 -12.045 ;
      RECT -1.805 -10.565 -1.705 -10.465 ;
      RECT -1.805 -10.325 -1.705 -10.225 ;
      RECT -1.805 -9.74 -1.705 -9.64 ;
      RECT -1.805 -0.05 -1.705 0.05 ;
      RECT -1.805 0.535 -1.705 0.635 ;
      RECT -1.805 0.775 -1.705 0.875 ;
      RECT -2.065 -55.905 -1.965 -55.805 ;
      RECT -2.065 -54.7 -1.965 -54.6 ;
      RECT -2.065 -51.145 -1.965 -51.045 ;
      RECT -2.065 -50.905 -1.965 -50.805 ;
      RECT -2.065 -49.325 -1.965 -49.225 ;
      RECT -2.065 -49.085 -1.965 -48.985 ;
      RECT -2.065 -45.53 -1.965 -45.43 ;
      RECT -2.065 -44.325 -1.965 -44.225 ;
      RECT -2.065 -42.985 -1.965 -42.885 ;
      RECT -2.065 -41.78 -1.965 -41.68 ;
      RECT -2.065 -38.225 -1.965 -38.125 ;
      RECT -2.065 -37.985 -1.965 -37.885 ;
      RECT -2.065 -36.405 -1.965 -36.305 ;
      RECT -2.065 -36.165 -1.965 -36.065 ;
      RECT -2.065 -32.61 -1.965 -32.51 ;
      RECT -2.065 -31.405 -1.965 -31.305 ;
      RECT -2.065 -30.065 -1.965 -29.965 ;
      RECT -2.065 -28.86 -1.965 -28.76 ;
      RECT -2.065 -25.305 -1.965 -25.205 ;
      RECT -2.065 -25.065 -1.965 -24.965 ;
      RECT -2.065 -23.485 -1.965 -23.385 ;
      RECT -2.065 -23.245 -1.965 -23.145 ;
      RECT -2.065 -19.69 -1.965 -19.59 ;
      RECT -2.065 -18.485 -1.965 -18.385 ;
      RECT -2.065 -17.145 -1.965 -17.045 ;
      RECT -2.065 -15.94 -1.965 -15.84 ;
      RECT -2.065 -12.385 -1.965 -12.285 ;
      RECT -2.065 -12.145 -1.965 -12.045 ;
      RECT -2.065 -10.565 -1.965 -10.465 ;
      RECT -2.065 -10.325 -1.965 -10.225 ;
      RECT -2.065 -6.77 -1.965 -6.67 ;
      RECT -2.065 -5.565 -1.965 -5.465 ;
      RECT -2.065 -4.225 -1.965 -4.125 ;
      RECT -2.065 -3.02 -1.965 -2.92 ;
      RECT -2.065 0.535 -1.965 0.635 ;
      RECT -2.065 0.775 -1.965 0.875 ;
      RECT -2.585 -55.905 -2.485 -55.805 ;
      RECT -2.585 -55.665 -2.485 -55.565 ;
      RECT -2.585 -51.73 -2.485 -51.63 ;
      RECT -2.585 -51.145 -2.485 -51.045 ;
      RECT -2.585 -50.905 -2.485 -50.805 ;
      RECT -2.585 -49.325 -2.485 -49.225 ;
      RECT -2.585 -49.085 -2.485 -48.985 ;
      RECT -2.585 -48.5 -2.485 -48.4 ;
      RECT -2.585 -44.565 -2.485 -44.465 ;
      RECT -2.585 -44.325 -2.485 -44.225 ;
      RECT -2.585 -42.985 -2.485 -42.885 ;
      RECT -2.585 -42.745 -2.485 -42.645 ;
      RECT -2.585 -38.81 -2.485 -38.71 ;
      RECT -2.585 -38.225 -2.485 -38.125 ;
      RECT -2.585 -37.985 -2.485 -37.885 ;
      RECT -2.585 -36.405 -2.485 -36.305 ;
      RECT -2.585 -36.165 -2.485 -36.065 ;
      RECT -2.585 -35.58 -2.485 -35.48 ;
      RECT -2.585 -31.645 -2.485 -31.545 ;
      RECT -2.585 -31.405 -2.485 -31.305 ;
      RECT -2.585 -30.065 -2.485 -29.965 ;
      RECT -2.585 -29.825 -2.485 -29.725 ;
      RECT -2.585 -25.89 -2.485 -25.79 ;
      RECT -2.585 -25.305 -2.485 -25.205 ;
      RECT -2.585 -25.065 -2.485 -24.965 ;
      RECT -2.585 -23.485 -2.485 -23.385 ;
      RECT -2.585 -23.245 -2.485 -23.145 ;
      RECT -2.585 -22.66 -2.485 -22.56 ;
      RECT -2.585 -18.725 -2.485 -18.625 ;
      RECT -2.585 -18.485 -2.485 -18.385 ;
      RECT -2.585 -17.145 -2.485 -17.045 ;
      RECT -2.585 -16.905 -2.485 -16.805 ;
      RECT -2.585 -12.97 -2.485 -12.87 ;
      RECT -2.585 -12.385 -2.485 -12.285 ;
      RECT -2.585 -12.145 -2.485 -12.045 ;
      RECT -2.585 -10.565 -2.485 -10.465 ;
      RECT -2.585 -10.325 -2.485 -10.225 ;
      RECT -2.585 -9.74 -2.485 -9.64 ;
      RECT -2.585 -5.805 -2.485 -5.705 ;
      RECT -2.585 -5.565 -2.485 -5.465 ;
      RECT -2.585 -4.225 -2.485 -4.125 ;
      RECT -2.585 -3.985 -2.485 -3.885 ;
      RECT -2.585 -0.05 -2.485 0.05 ;
      RECT -2.585 0.535 -2.485 0.635 ;
      RECT -2.585 0.775 -2.485 0.875 ;
      RECT -3.105 -51.73 -3.005 -51.63 ;
      RECT -3.105 -51.145 -3.005 -51.045 ;
      RECT -3.105 -50.905 -3.005 -50.805 ;
      RECT -3.105 -49.325 -3.005 -49.225 ;
      RECT -3.105 -49.085 -3.005 -48.985 ;
      RECT -3.105 -48.5 -3.005 -48.4 ;
      RECT -3.105 -38.81 -3.005 -38.71 ;
      RECT -3.105 -38.225 -3.005 -38.125 ;
      RECT -3.105 -37.985 -3.005 -37.885 ;
      RECT -3.105 -36.405 -3.005 -36.305 ;
      RECT -3.105 -36.165 -3.005 -36.065 ;
      RECT -3.105 -35.58 -3.005 -35.48 ;
      RECT -3.105 -25.89 -3.005 -25.79 ;
      RECT -3.105 -25.305 -3.005 -25.205 ;
      RECT -3.105 -25.065 -3.005 -24.965 ;
      RECT -3.105 -23.485 -3.005 -23.385 ;
      RECT -3.105 -23.245 -3.005 -23.145 ;
      RECT -3.105 -22.66 -3.005 -22.56 ;
      RECT -3.105 -12.97 -3.005 -12.87 ;
      RECT -3.105 -12.385 -3.005 -12.285 ;
      RECT -3.105 -12.145 -3.005 -12.045 ;
      RECT -3.105 -10.565 -3.005 -10.465 ;
      RECT -3.105 -10.325 -3.005 -10.225 ;
      RECT -3.105 -9.74 -3.005 -9.64 ;
      RECT -3.105 -0.05 -3.005 0.05 ;
      RECT -3.105 0.535 -3.005 0.635 ;
      RECT -3.105 0.775 -3.005 0.875 ;
      RECT -3.365 -55.905 -3.265 -55.805 ;
      RECT -3.365 -51.99 -3.265 -51.89 ;
      RECT -3.365 -51.145 -3.265 -51.045 ;
      RECT -3.365 -50.905 -3.265 -50.805 ;
      RECT -3.365 -49.325 -3.265 -49.225 ;
      RECT -3.365 -49.085 -3.265 -48.985 ;
      RECT -3.365 -48.24 -3.265 -48.14 ;
      RECT -3.365 -44.325 -3.265 -44.225 ;
      RECT -3.365 -42.985 -3.265 -42.885 ;
      RECT -3.365 -39.07 -3.265 -38.97 ;
      RECT -3.365 -38.225 -3.265 -38.125 ;
      RECT -3.365 -37.985 -3.265 -37.885 ;
      RECT -3.365 -36.405 -3.265 -36.305 ;
      RECT -3.365 -36.165 -3.265 -36.065 ;
      RECT -3.365 -35.32 -3.265 -35.22 ;
      RECT -3.365 -31.405 -3.265 -31.305 ;
      RECT -3.365 -30.065 -3.265 -29.965 ;
      RECT -3.365 -26.15 -3.265 -26.05 ;
      RECT -3.365 -25.305 -3.265 -25.205 ;
      RECT -3.365 -25.065 -3.265 -24.965 ;
      RECT -3.365 -23.485 -3.265 -23.385 ;
      RECT -3.365 -23.245 -3.265 -23.145 ;
      RECT -3.365 -22.4 -3.265 -22.3 ;
      RECT -3.365 -18.485 -3.265 -18.385 ;
      RECT -3.365 -17.145 -3.265 -17.045 ;
      RECT -3.365 -13.23 -3.265 -13.13 ;
      RECT -3.365 -12.385 -3.265 -12.285 ;
      RECT -3.365 -12.145 -3.265 -12.045 ;
      RECT -3.365 -10.565 -3.265 -10.465 ;
      RECT -3.365 -10.325 -3.265 -10.225 ;
      RECT -3.365 -9.48 -3.265 -9.38 ;
      RECT -3.365 -5.565 -3.265 -5.465 ;
      RECT -3.365 -4.225 -3.265 -4.125 ;
      RECT -3.365 -0.31 -3.265 -0.21 ;
      RECT -3.365 0.535 -3.265 0.635 ;
      RECT -3.365 0.775 -3.265 0.875 ;
      RECT -3.885 -55.905 -3.785 -55.805 ;
      RECT -3.885 -55.665 -3.785 -55.565 ;
      RECT -3.885 -51.73 -3.785 -51.63 ;
      RECT -3.885 -51.145 -3.785 -51.045 ;
      RECT -3.885 -50.905 -3.785 -50.805 ;
      RECT -3.885 -49.325 -3.785 -49.225 ;
      RECT -3.885 -49.085 -3.785 -48.985 ;
      RECT -3.885 -48.5 -3.785 -48.4 ;
      RECT -3.885 -44.565 -3.785 -44.465 ;
      RECT -3.885 -44.325 -3.785 -44.225 ;
      RECT -3.885 -42.985 -3.785 -42.885 ;
      RECT -3.885 -42.745 -3.785 -42.645 ;
      RECT -3.885 -38.81 -3.785 -38.71 ;
      RECT -3.885 -38.225 -3.785 -38.125 ;
      RECT -3.885 -37.985 -3.785 -37.885 ;
      RECT -3.885 -36.405 -3.785 -36.305 ;
      RECT -3.885 -36.165 -3.785 -36.065 ;
      RECT -3.885 -35.58 -3.785 -35.48 ;
      RECT -3.885 -31.645 -3.785 -31.545 ;
      RECT -3.885 -31.405 -3.785 -31.305 ;
      RECT -3.885 -30.065 -3.785 -29.965 ;
      RECT -3.885 -29.825 -3.785 -29.725 ;
      RECT -3.885 -25.89 -3.785 -25.79 ;
      RECT -3.885 -25.305 -3.785 -25.205 ;
      RECT -3.885 -25.065 -3.785 -24.965 ;
      RECT -3.885 -23.485 -3.785 -23.385 ;
      RECT -3.885 -23.245 -3.785 -23.145 ;
      RECT -3.885 -22.66 -3.785 -22.56 ;
      RECT -3.885 -18.725 -3.785 -18.625 ;
      RECT -3.885 -18.485 -3.785 -18.385 ;
      RECT -3.885 -17.145 -3.785 -17.045 ;
      RECT -3.885 -16.905 -3.785 -16.805 ;
      RECT -3.885 -12.97 -3.785 -12.87 ;
      RECT -3.885 -12.385 -3.785 -12.285 ;
      RECT -3.885 -12.145 -3.785 -12.045 ;
      RECT -3.885 -10.565 -3.785 -10.465 ;
      RECT -3.885 -10.325 -3.785 -10.225 ;
      RECT -3.885 -9.74 -3.785 -9.64 ;
      RECT -3.885 -5.805 -3.785 -5.705 ;
      RECT -3.885 -5.565 -3.785 -5.465 ;
      RECT -3.885 -4.225 -3.785 -4.125 ;
      RECT -3.885 -3.985 -3.785 -3.885 ;
      RECT -3.885 -0.05 -3.785 0.05 ;
      RECT -3.885 0.535 -3.785 0.635 ;
      RECT -3.885 0.775 -3.785 0.875 ;
      RECT -4.405 -51.73 -4.305 -51.63 ;
      RECT -4.405 -51.145 -4.305 -51.045 ;
      RECT -4.405 -50.905 -4.305 -50.805 ;
      RECT -4.405 -49.325 -4.305 -49.225 ;
      RECT -4.405 -49.085 -4.305 -48.985 ;
      RECT -4.405 -48.5 -4.305 -48.4 ;
      RECT -4.405 -38.81 -4.305 -38.71 ;
      RECT -4.405 -38.225 -4.305 -38.125 ;
      RECT -4.405 -37.985 -4.305 -37.885 ;
      RECT -4.405 -36.405 -4.305 -36.305 ;
      RECT -4.405 -36.165 -4.305 -36.065 ;
      RECT -4.405 -35.58 -4.305 -35.48 ;
      RECT -4.405 -25.89 -4.305 -25.79 ;
      RECT -4.405 -25.305 -4.305 -25.205 ;
      RECT -4.405 -25.065 -4.305 -24.965 ;
      RECT -4.405 -23.485 -4.305 -23.385 ;
      RECT -4.405 -23.245 -4.305 -23.145 ;
      RECT -4.405 -22.66 -4.305 -22.56 ;
      RECT -4.405 -12.97 -4.305 -12.87 ;
      RECT -4.405 -12.385 -4.305 -12.285 ;
      RECT -4.405 -12.145 -4.305 -12.045 ;
      RECT -4.405 -10.565 -4.305 -10.465 ;
      RECT -4.405 -10.325 -4.305 -10.225 ;
      RECT -4.405 -9.74 -4.305 -9.64 ;
      RECT -4.405 -0.05 -4.305 0.05 ;
      RECT -4.405 0.535 -4.305 0.635 ;
      RECT -4.405 0.775 -4.305 0.875 ;
      RECT -4.665 -55.905 -4.565 -55.805 ;
      RECT -4.665 -51.47 -4.565 -51.37 ;
      RECT -4.665 -51.145 -4.565 -51.045 ;
      RECT -4.665 -50.905 -4.565 -50.805 ;
      RECT -4.665 -49.325 -4.565 -49.225 ;
      RECT -4.665 -49.085 -4.565 -48.985 ;
      RECT -4.665 -48.76 -4.565 -48.66 ;
      RECT -4.665 -44.325 -4.565 -44.225 ;
      RECT -4.665 -42.985 -4.565 -42.885 ;
      RECT -4.665 -38.55 -4.565 -38.45 ;
      RECT -4.665 -38.225 -4.565 -38.125 ;
      RECT -4.665 -37.985 -4.565 -37.885 ;
      RECT -4.665 -36.405 -4.565 -36.305 ;
      RECT -4.665 -36.165 -4.565 -36.065 ;
      RECT -4.665 -35.84 -4.565 -35.74 ;
      RECT -4.665 -31.405 -4.565 -31.305 ;
      RECT -4.665 -30.065 -4.565 -29.965 ;
      RECT -4.665 -25.63 -4.565 -25.53 ;
      RECT -4.665 -25.305 -4.565 -25.205 ;
      RECT -4.665 -25.065 -4.565 -24.965 ;
      RECT -4.665 -23.485 -4.565 -23.385 ;
      RECT -4.665 -23.245 -4.565 -23.145 ;
      RECT -4.665 -22.92 -4.565 -22.82 ;
      RECT -4.665 -18.485 -4.565 -18.385 ;
      RECT -4.665 -17.145 -4.565 -17.045 ;
      RECT -4.665 -12.71 -4.565 -12.61 ;
      RECT -4.665 -12.385 -4.565 -12.285 ;
      RECT -4.665 -12.145 -4.565 -12.045 ;
      RECT -4.665 -10.565 -4.565 -10.465 ;
      RECT -4.665 -10.325 -4.565 -10.225 ;
      RECT -4.665 -10 -4.565 -9.9 ;
      RECT -4.665 -5.565 -4.565 -5.465 ;
      RECT -4.665 -4.225 -4.565 -4.125 ;
      RECT -4.665 0.21 -4.565 0.31 ;
      RECT -4.665 0.535 -4.565 0.635 ;
      RECT -4.665 0.775 -4.565 0.875 ;
      RECT -4.925 -59.27 -4.825 -59.17 ;
      RECT -4.925 -52.315 -4.825 -52.215 ;
      RECT -4.925 -47.695 -4.825 -47.595 ;
      RECT -4.925 -39.615 -4.825 -39.515 ;
      RECT -4.925 -34.775 -4.825 -34.675 ;
      RECT -4.925 -26.695 -4.825 -26.595 ;
      RECT -4.925 -21.855 -4.825 -21.755 ;
      RECT -4.925 -13.775 -4.825 -13.675 ;
      RECT -4.925 -8.935 -4.825 -8.835 ;
      RECT -4.925 -0.855 -4.825 -0.755 ;
      RECT -4.925 4.135 -4.825 4.235 ;
      RECT -5.185 -55.905 -5.085 -55.805 ;
      RECT -5.185 -55.665 -5.085 -55.565 ;
      RECT -5.185 -51.73 -5.085 -51.63 ;
      RECT -5.185 -51.145 -5.085 -51.045 ;
      RECT -5.185 -50.905 -5.085 -50.805 ;
      RECT -5.185 -49.325 -5.085 -49.225 ;
      RECT -5.185 -49.085 -5.085 -48.985 ;
      RECT -5.185 -48.5 -5.085 -48.4 ;
      RECT -5.185 -44.565 -5.085 -44.465 ;
      RECT -5.185 -44.325 -5.085 -44.225 ;
      RECT -5.185 -42.985 -5.085 -42.885 ;
      RECT -5.185 -42.745 -5.085 -42.645 ;
      RECT -5.185 -38.81 -5.085 -38.71 ;
      RECT -5.185 -38.225 -5.085 -38.125 ;
      RECT -5.185 -37.985 -5.085 -37.885 ;
      RECT -5.185 -36.405 -5.085 -36.305 ;
      RECT -5.185 -36.165 -5.085 -36.065 ;
      RECT -5.185 -35.58 -5.085 -35.48 ;
      RECT -5.185 -31.645 -5.085 -31.545 ;
      RECT -5.185 -31.405 -5.085 -31.305 ;
      RECT -5.185 -30.065 -5.085 -29.965 ;
      RECT -5.185 -29.825 -5.085 -29.725 ;
      RECT -5.185 -25.89 -5.085 -25.79 ;
      RECT -5.185 -25.305 -5.085 -25.205 ;
      RECT -5.185 -25.065 -5.085 -24.965 ;
      RECT -5.185 -23.485 -5.085 -23.385 ;
      RECT -5.185 -23.245 -5.085 -23.145 ;
      RECT -5.185 -22.66 -5.085 -22.56 ;
      RECT -5.185 -18.725 -5.085 -18.625 ;
      RECT -5.185 -18.485 -5.085 -18.385 ;
      RECT -5.185 -17.145 -5.085 -17.045 ;
      RECT -5.185 -16.905 -5.085 -16.805 ;
      RECT -5.185 -12.97 -5.085 -12.87 ;
      RECT -5.185 -12.385 -5.085 -12.285 ;
      RECT -5.185 -12.145 -5.085 -12.045 ;
      RECT -5.185 -10.565 -5.085 -10.465 ;
      RECT -5.185 -10.325 -5.085 -10.225 ;
      RECT -5.185 -9.74 -5.085 -9.64 ;
      RECT -5.185 -5.805 -5.085 -5.705 ;
      RECT -5.185 -5.565 -5.085 -5.465 ;
      RECT -5.185 -4.225 -5.085 -4.125 ;
      RECT -5.185 -3.985 -5.085 -3.885 ;
      RECT -5.185 -0.05 -5.085 0.05 ;
      RECT -5.185 0.535 -5.085 0.635 ;
      RECT -5.185 0.775 -5.085 0.875 ;
      RECT -5.705 -51.73 -5.605 -51.63 ;
      RECT -5.705 -51.145 -5.605 -51.045 ;
      RECT -5.705 -50.905 -5.605 -50.805 ;
      RECT -5.705 -49.325 -5.605 -49.225 ;
      RECT -5.705 -49.085 -5.605 -48.985 ;
      RECT -5.705 -48.5 -5.605 -48.4 ;
      RECT -5.705 -38.81 -5.605 -38.71 ;
      RECT -5.705 -38.225 -5.605 -38.125 ;
      RECT -5.705 -37.985 -5.605 -37.885 ;
      RECT -5.705 -36.405 -5.605 -36.305 ;
      RECT -5.705 -36.165 -5.605 -36.065 ;
      RECT -5.705 -35.58 -5.605 -35.48 ;
      RECT -5.705 -25.89 -5.605 -25.79 ;
      RECT -5.705 -25.305 -5.605 -25.205 ;
      RECT -5.705 -25.065 -5.605 -24.965 ;
      RECT -5.705 -23.485 -5.605 -23.385 ;
      RECT -5.705 -23.245 -5.605 -23.145 ;
      RECT -5.705 -22.66 -5.605 -22.56 ;
      RECT -5.705 -12.97 -5.605 -12.87 ;
      RECT -5.705 -12.385 -5.605 -12.285 ;
      RECT -5.705 -12.145 -5.605 -12.045 ;
      RECT -5.705 -10.565 -5.605 -10.465 ;
      RECT -5.705 -10.325 -5.605 -10.225 ;
      RECT -5.705 -9.74 -5.605 -9.64 ;
      RECT -5.705 -0.05 -5.605 0.05 ;
      RECT -5.705 0.535 -5.605 0.635 ;
      RECT -5.705 0.775 -5.605 0.875 ;
      RECT -5.965 -55.905 -5.865 -55.805 ;
      RECT -5.965 -52.535 -5.865 -52.435 ;
      RECT -5.965 -51.145 -5.865 -51.045 ;
      RECT -5.965 -50.905 -5.865 -50.805 ;
      RECT -5.965 -49.325 -5.865 -49.225 ;
      RECT -5.965 -49.085 -5.865 -48.985 ;
      RECT -5.965 -46.815 -5.865 -46.715 ;
      RECT -5.965 -44.325 -5.865 -44.225 ;
      RECT -5.965 -42.985 -5.865 -42.885 ;
      RECT -5.965 -40.495 -5.865 -40.395 ;
      RECT -5.965 -38.225 -5.865 -38.125 ;
      RECT -5.965 -37.985 -5.865 -37.885 ;
      RECT -5.965 -36.405 -5.865 -36.305 ;
      RECT -5.965 -36.165 -5.865 -36.065 ;
      RECT -5.965 -33.895 -5.865 -33.795 ;
      RECT -5.965 -31.405 -5.865 -31.305 ;
      RECT -5.965 -30.065 -5.865 -29.965 ;
      RECT -5.965 -27.575 -5.865 -27.475 ;
      RECT -5.965 -25.305 -5.865 -25.205 ;
      RECT -5.965 -25.065 -5.865 -24.965 ;
      RECT -5.965 -23.485 -5.865 -23.385 ;
      RECT -5.965 -23.245 -5.865 -23.145 ;
      RECT -5.965 -20.975 -5.865 -20.875 ;
      RECT -5.965 -18.485 -5.865 -18.385 ;
      RECT -5.965 -17.145 -5.865 -17.045 ;
      RECT -5.965 -14.655 -5.865 -14.555 ;
      RECT -5.965 -12.385 -5.865 -12.285 ;
      RECT -5.965 -12.145 -5.865 -12.045 ;
      RECT -5.965 -10.565 -5.865 -10.465 ;
      RECT -5.965 -10.325 -5.865 -10.225 ;
      RECT -5.965 -8.055 -5.865 -7.955 ;
      RECT -5.965 -5.565 -5.865 -5.465 ;
      RECT -5.965 -4.225 -5.865 -4.125 ;
      RECT -5.965 -1.735 -5.865 -1.635 ;
      RECT -5.965 0.535 -5.865 0.635 ;
      RECT -5.965 0.775 -5.865 0.875 ;
      RECT -6.485 -55.905 -6.385 -55.805 ;
      RECT -6.485 -55.665 -6.385 -55.565 ;
      RECT -6.485 -51.435 -6.385 -51.335 ;
      RECT -6.485 -51.145 -6.385 -51.045 ;
      RECT -6.485 -50.905 -6.385 -50.805 ;
      RECT -6.485 -49.325 -6.385 -49.225 ;
      RECT -6.485 -49.085 -6.385 -48.985 ;
      RECT -6.485 -48.795 -6.385 -48.695 ;
      RECT -6.485 -44.565 -6.385 -44.465 ;
      RECT -6.485 -44.325 -6.385 -44.225 ;
      RECT -6.485 -42.985 -6.385 -42.885 ;
      RECT -6.485 -42.745 -6.385 -42.645 ;
      RECT -6.485 -38.515 -6.385 -38.415 ;
      RECT -6.485 -38.225 -6.385 -38.125 ;
      RECT -6.485 -37.985 -6.385 -37.885 ;
      RECT -6.485 -36.405 -6.385 -36.305 ;
      RECT -6.485 -36.165 -6.385 -36.065 ;
      RECT -6.485 -35.875 -6.385 -35.775 ;
      RECT -6.485 -31.645 -6.385 -31.545 ;
      RECT -6.485 -31.405 -6.385 -31.305 ;
      RECT -6.485 -30.065 -6.385 -29.965 ;
      RECT -6.485 -29.825 -6.385 -29.725 ;
      RECT -6.485 -25.595 -6.385 -25.495 ;
      RECT -6.485 -25.305 -6.385 -25.205 ;
      RECT -6.485 -25.065 -6.385 -24.965 ;
      RECT -6.485 -23.485 -6.385 -23.385 ;
      RECT -6.485 -23.245 -6.385 -23.145 ;
      RECT -6.485 -22.955 -6.385 -22.855 ;
      RECT -6.485 -18.725 -6.385 -18.625 ;
      RECT -6.485 -18.485 -6.385 -18.385 ;
      RECT -6.485 -17.145 -6.385 -17.045 ;
      RECT -6.485 -16.905 -6.385 -16.805 ;
      RECT -6.485 -12.675 -6.385 -12.575 ;
      RECT -6.485 -12.385 -6.385 -12.285 ;
      RECT -6.485 -12.145 -6.385 -12.045 ;
      RECT -6.485 -10.565 -6.385 -10.465 ;
      RECT -6.485 -10.325 -6.385 -10.225 ;
      RECT -6.485 -10.035 -6.385 -9.935 ;
      RECT -6.485 -5.805 -6.385 -5.705 ;
      RECT -6.485 -5.565 -6.385 -5.465 ;
      RECT -6.485 -4.225 -6.385 -4.125 ;
      RECT -6.485 -3.985 -6.385 -3.885 ;
      RECT -6.485 0.245 -6.385 0.345 ;
      RECT -6.485 0.535 -6.385 0.635 ;
      RECT -6.485 0.775 -6.385 0.875 ;
      RECT -7.265 -55.905 -7.165 -55.805 ;
      RECT -7.265 -52.095 -7.165 -51.995 ;
      RECT -7.265 -51.145 -7.165 -51.045 ;
      RECT -7.265 -50.905 -7.165 -50.805 ;
      RECT -7.265 -49.325 -7.165 -49.225 ;
      RECT -7.265 -49.085 -7.165 -48.985 ;
      RECT -7.265 -47.035 -7.165 -46.935 ;
      RECT -7.265 -44.325 -7.165 -44.225 ;
      RECT -7.265 -42.985 -7.165 -42.885 ;
      RECT -7.265 -40.275 -7.165 -40.175 ;
      RECT -7.265 -38.225 -7.165 -38.125 ;
      RECT -7.265 -37.985 -7.165 -37.885 ;
      RECT -7.265 -36.405 -7.165 -36.305 ;
      RECT -7.265 -36.165 -7.165 -36.065 ;
      RECT -7.265 -34.115 -7.165 -34.015 ;
      RECT -7.265 -31.405 -7.165 -31.305 ;
      RECT -7.265 -30.065 -7.165 -29.965 ;
      RECT -7.265 -27.355 -7.165 -27.255 ;
      RECT -7.265 -25.305 -7.165 -25.205 ;
      RECT -7.265 -25.065 -7.165 -24.965 ;
      RECT -7.265 -23.485 -7.165 -23.385 ;
      RECT -7.265 -23.245 -7.165 -23.145 ;
      RECT -7.265 -21.195 -7.165 -21.095 ;
      RECT -7.265 -18.485 -7.165 -18.385 ;
      RECT -7.265 -17.145 -7.165 -17.045 ;
      RECT -7.265 -14.435 -7.165 -14.335 ;
      RECT -7.265 -12.385 -7.165 -12.285 ;
      RECT -7.265 -12.145 -7.165 -12.045 ;
      RECT -7.265 -10.565 -7.165 -10.465 ;
      RECT -7.265 -10.325 -7.165 -10.225 ;
      RECT -7.265 -8.275 -7.165 -8.175 ;
      RECT -7.265 -5.565 -7.165 -5.465 ;
      RECT -7.265 -4.225 -7.165 -4.125 ;
      RECT -7.265 -1.515 -7.165 -1.415 ;
      RECT -7.265 0.535 -7.165 0.635 ;
      RECT -7.265 0.775 -7.165 0.875 ;
      RECT -7.785 -55.905 -7.685 -55.805 ;
      RECT -7.785 -55.665 -7.685 -55.565 ;
      RECT -7.785 -51.435 -7.685 -51.335 ;
      RECT -7.785 -51.145 -7.685 -51.045 ;
      RECT -7.785 -50.905 -7.685 -50.805 ;
      RECT -7.785 -49.325 -7.685 -49.225 ;
      RECT -7.785 -49.085 -7.685 -48.985 ;
      RECT -7.785 -48.795 -7.685 -48.695 ;
      RECT -7.785 -44.565 -7.685 -44.465 ;
      RECT -7.785 -44.325 -7.685 -44.225 ;
      RECT -7.785 -42.985 -7.685 -42.885 ;
      RECT -7.785 -42.745 -7.685 -42.645 ;
      RECT -7.785 -38.515 -7.685 -38.415 ;
      RECT -7.785 -38.225 -7.685 -38.125 ;
      RECT -7.785 -37.985 -7.685 -37.885 ;
      RECT -7.785 -36.405 -7.685 -36.305 ;
      RECT -7.785 -36.165 -7.685 -36.065 ;
      RECT -7.785 -35.875 -7.685 -35.775 ;
      RECT -7.785 -31.645 -7.685 -31.545 ;
      RECT -7.785 -31.405 -7.685 -31.305 ;
      RECT -7.785 -30.065 -7.685 -29.965 ;
      RECT -7.785 -29.825 -7.685 -29.725 ;
      RECT -7.785 -25.595 -7.685 -25.495 ;
      RECT -7.785 -25.305 -7.685 -25.205 ;
      RECT -7.785 -25.065 -7.685 -24.965 ;
      RECT -7.785 -23.485 -7.685 -23.385 ;
      RECT -7.785 -23.245 -7.685 -23.145 ;
      RECT -7.785 -22.955 -7.685 -22.855 ;
      RECT -7.785 -18.725 -7.685 -18.625 ;
      RECT -7.785 -18.485 -7.685 -18.385 ;
      RECT -7.785 -17.145 -7.685 -17.045 ;
      RECT -7.785 -16.905 -7.685 -16.805 ;
      RECT -7.785 -12.675 -7.685 -12.575 ;
      RECT -7.785 -12.385 -7.685 -12.285 ;
      RECT -7.785 -12.145 -7.685 -12.045 ;
      RECT -7.785 -10.565 -7.685 -10.465 ;
      RECT -7.785 -10.325 -7.685 -10.225 ;
      RECT -7.785 -10.035 -7.685 -9.935 ;
      RECT -7.785 -5.805 -7.685 -5.705 ;
      RECT -7.785 -5.565 -7.685 -5.465 ;
      RECT -7.785 -4.225 -7.685 -4.125 ;
      RECT -7.785 -3.985 -7.685 -3.885 ;
      RECT -7.785 0.245 -7.685 0.345 ;
      RECT -7.785 0.535 -7.685 0.635 ;
      RECT -7.785 0.775 -7.685 0.875 ;
      RECT -8.565 -55.905 -8.465 -55.805 ;
      RECT -8.565 -52.975 -8.465 -52.875 ;
      RECT -8.565 -51.145 -8.465 -51.045 ;
      RECT -8.565 -50.905 -8.465 -50.805 ;
      RECT -8.565 -49.325 -8.465 -49.225 ;
      RECT -8.565 -49.085 -8.465 -48.985 ;
      RECT -8.565 -46.815 -8.465 -46.715 ;
      RECT -8.565 -44.325 -8.465 -44.225 ;
      RECT -8.565 -42.985 -8.465 -42.885 ;
      RECT -8.565 -40.495 -8.465 -40.395 ;
      RECT -8.565 -38.225 -8.465 -38.125 ;
      RECT -8.565 -37.985 -8.465 -37.885 ;
      RECT -8.565 -36.405 -8.465 -36.305 ;
      RECT -8.565 -36.165 -8.465 -36.065 ;
      RECT -8.565 -33.895 -8.465 -33.795 ;
      RECT -8.565 -31.405 -8.465 -31.305 ;
      RECT -8.565 -30.065 -8.465 -29.965 ;
      RECT -8.565 -27.575 -8.465 -27.475 ;
      RECT -8.565 -25.305 -8.465 -25.205 ;
      RECT -8.565 -25.065 -8.465 -24.965 ;
      RECT -8.565 -23.485 -8.465 -23.385 ;
      RECT -8.565 -23.245 -8.465 -23.145 ;
      RECT -8.565 -20.975 -8.465 -20.875 ;
      RECT -8.565 -18.485 -8.465 -18.385 ;
      RECT -8.565 -17.145 -8.465 -17.045 ;
      RECT -8.565 -14.655 -8.465 -14.555 ;
      RECT -8.565 -12.385 -8.465 -12.285 ;
      RECT -8.565 -12.145 -8.465 -12.045 ;
      RECT -8.565 -10.565 -8.465 -10.465 ;
      RECT -8.565 -10.325 -8.465 -10.225 ;
      RECT -8.565 -8.055 -8.465 -7.955 ;
      RECT -8.565 -5.565 -8.465 -5.465 ;
      RECT -8.565 -4.225 -8.465 -4.125 ;
      RECT -8.565 -1.735 -8.465 -1.635 ;
      RECT -8.565 0.535 -8.465 0.635 ;
      RECT -8.565 0.775 -8.465 0.875 ;
      RECT -9.085 -55.905 -8.985 -55.805 ;
      RECT -9.085 -55.665 -8.985 -55.565 ;
      RECT -9.085 -51.435 -8.985 -51.335 ;
      RECT -9.085 -51.145 -8.985 -51.045 ;
      RECT -9.085 -50.905 -8.985 -50.805 ;
      RECT -9.085 -49.325 -8.985 -49.225 ;
      RECT -9.085 -49.085 -8.985 -48.985 ;
      RECT -9.085 -48.795 -8.985 -48.695 ;
      RECT -9.085 -44.565 -8.985 -44.465 ;
      RECT -9.085 -44.325 -8.985 -44.225 ;
      RECT -9.085 -42.985 -8.985 -42.885 ;
      RECT -9.085 -42.745 -8.985 -42.645 ;
      RECT -9.085 -38.515 -8.985 -38.415 ;
      RECT -9.085 -38.225 -8.985 -38.125 ;
      RECT -9.085 -37.985 -8.985 -37.885 ;
      RECT -9.085 -36.405 -8.985 -36.305 ;
      RECT -9.085 -36.165 -8.985 -36.065 ;
      RECT -9.085 -35.875 -8.985 -35.775 ;
      RECT -9.085 -31.645 -8.985 -31.545 ;
      RECT -9.085 -31.405 -8.985 -31.305 ;
      RECT -9.085 -30.065 -8.985 -29.965 ;
      RECT -9.085 -29.825 -8.985 -29.725 ;
      RECT -9.085 -25.595 -8.985 -25.495 ;
      RECT -9.085 -25.305 -8.985 -25.205 ;
      RECT -9.085 -25.065 -8.985 -24.965 ;
      RECT -9.085 -23.485 -8.985 -23.385 ;
      RECT -9.085 -23.245 -8.985 -23.145 ;
      RECT -9.085 -22.955 -8.985 -22.855 ;
      RECT -9.085 -18.725 -8.985 -18.625 ;
      RECT -9.085 -18.485 -8.985 -18.385 ;
      RECT -9.085 -17.145 -8.985 -17.045 ;
      RECT -9.085 -16.905 -8.985 -16.805 ;
      RECT -9.085 -12.675 -8.985 -12.575 ;
      RECT -9.085 -12.385 -8.985 -12.285 ;
      RECT -9.085 -12.145 -8.985 -12.045 ;
      RECT -9.085 -10.565 -8.985 -10.465 ;
      RECT -9.085 -10.325 -8.985 -10.225 ;
      RECT -9.085 -10.035 -8.985 -9.935 ;
      RECT -9.085 -5.805 -8.985 -5.705 ;
      RECT -9.085 -5.565 -8.985 -5.465 ;
      RECT -9.085 -4.225 -8.985 -4.125 ;
      RECT -9.085 -3.985 -8.985 -3.885 ;
      RECT -9.085 0.245 -8.985 0.345 ;
      RECT -9.085 0.535 -8.985 0.635 ;
      RECT -9.085 0.775 -8.985 0.875 ;
      RECT -9.865 -55.905 -9.765 -55.805 ;
      RECT -9.865 -52.755 -9.765 -52.655 ;
      RECT -9.865 -51.145 -9.765 -51.045 ;
      RECT -9.865 -50.905 -9.765 -50.805 ;
      RECT -9.865 -49.325 -9.765 -49.225 ;
      RECT -9.865 -49.085 -9.765 -48.985 ;
      RECT -9.865 -47.035 -9.765 -46.935 ;
      RECT -9.865 -44.325 -9.765 -44.225 ;
      RECT -9.865 -42.985 -9.765 -42.885 ;
      RECT -9.865 -40.275 -9.765 -40.175 ;
      RECT -9.865 -38.225 -9.765 -38.125 ;
      RECT -9.865 -37.985 -9.765 -37.885 ;
      RECT -9.865 -36.405 -9.765 -36.305 ;
      RECT -9.865 -36.165 -9.765 -36.065 ;
      RECT -9.865 -34.115 -9.765 -34.015 ;
      RECT -9.865 -31.405 -9.765 -31.305 ;
      RECT -9.865 -30.065 -9.765 -29.965 ;
      RECT -9.865 -27.355 -9.765 -27.255 ;
      RECT -9.865 -25.305 -9.765 -25.205 ;
      RECT -9.865 -25.065 -9.765 -24.965 ;
      RECT -9.865 -23.485 -9.765 -23.385 ;
      RECT -9.865 -23.245 -9.765 -23.145 ;
      RECT -9.865 -21.195 -9.765 -21.095 ;
      RECT -9.865 -18.485 -9.765 -18.385 ;
      RECT -9.865 -17.145 -9.765 -17.045 ;
      RECT -9.865 -14.435 -9.765 -14.335 ;
      RECT -9.865 -12.385 -9.765 -12.285 ;
      RECT -9.865 -12.145 -9.765 -12.045 ;
      RECT -9.865 -10.565 -9.765 -10.465 ;
      RECT -9.865 -10.325 -9.765 -10.225 ;
      RECT -9.865 -8.275 -9.765 -8.175 ;
      RECT -9.865 -5.565 -9.765 -5.465 ;
      RECT -9.865 -4.225 -9.765 -4.125 ;
      RECT -9.865 -1.515 -9.765 -1.415 ;
      RECT -9.865 0.535 -9.765 0.635 ;
      RECT -9.865 0.775 -9.765 0.875 ;
      RECT -10.385 -55.905 -10.285 -55.805 ;
      RECT -10.385 -55.665 -10.285 -55.565 ;
      RECT -10.385 -51.435 -10.285 -51.335 ;
      RECT -10.385 -51.145 -10.285 -51.045 ;
      RECT -10.385 -50.905 -10.285 -50.805 ;
      RECT -10.385 -49.325 -10.285 -49.225 ;
      RECT -10.385 -49.085 -10.285 -48.985 ;
      RECT -10.385 -48.795 -10.285 -48.695 ;
      RECT -10.385 -44.565 -10.285 -44.465 ;
      RECT -10.385 -44.325 -10.285 -44.225 ;
      RECT -10.385 -42.985 -10.285 -42.885 ;
      RECT -10.385 -42.745 -10.285 -42.645 ;
      RECT -10.385 -38.515 -10.285 -38.415 ;
      RECT -10.385 -38.225 -10.285 -38.125 ;
      RECT -10.385 -37.985 -10.285 -37.885 ;
      RECT -10.385 -36.405 -10.285 -36.305 ;
      RECT -10.385 -36.165 -10.285 -36.065 ;
      RECT -10.385 -35.875 -10.285 -35.775 ;
      RECT -10.385 -31.645 -10.285 -31.545 ;
      RECT -10.385 -31.405 -10.285 -31.305 ;
      RECT -10.385 -30.065 -10.285 -29.965 ;
      RECT -10.385 -29.825 -10.285 -29.725 ;
      RECT -10.385 -25.595 -10.285 -25.495 ;
      RECT -10.385 -25.305 -10.285 -25.205 ;
      RECT -10.385 -25.065 -10.285 -24.965 ;
      RECT -10.385 -23.485 -10.285 -23.385 ;
      RECT -10.385 -23.245 -10.285 -23.145 ;
      RECT -10.385 -22.955 -10.285 -22.855 ;
      RECT -10.385 -18.725 -10.285 -18.625 ;
      RECT -10.385 -18.485 -10.285 -18.385 ;
      RECT -10.385 -17.145 -10.285 -17.045 ;
      RECT -10.385 -16.905 -10.285 -16.805 ;
      RECT -10.385 -12.675 -10.285 -12.575 ;
      RECT -10.385 -12.385 -10.285 -12.285 ;
      RECT -10.385 -12.145 -10.285 -12.045 ;
      RECT -10.385 -10.565 -10.285 -10.465 ;
      RECT -10.385 -10.325 -10.285 -10.225 ;
      RECT -10.385 -10.035 -10.285 -9.935 ;
      RECT -10.385 -5.805 -10.285 -5.705 ;
      RECT -10.385 -5.565 -10.285 -5.465 ;
      RECT -10.385 -4.225 -10.285 -4.125 ;
      RECT -10.385 -3.985 -10.285 -3.885 ;
      RECT -10.385 0.245 -10.285 0.345 ;
      RECT -10.385 0.535 -10.285 0.635 ;
      RECT -10.385 0.775 -10.285 0.875 ;
      RECT -11.165 -49.325 -11.065 -49.225 ;
      RECT -11.165 -49.085 -11.065 -48.985 ;
      RECT -11.165 -48.135 -11.065 -48.035 ;
      RECT -11.165 -44.325 -11.065 -44.225 ;
      RECT -11.165 -42.985 -11.065 -42.885 ;
      RECT -11.165 -39.175 -11.065 -39.075 ;
      RECT -11.165 -38.225 -11.065 -38.125 ;
      RECT -11.165 -37.985 -11.065 -37.885 ;
      RECT -11.165 -36.405 -11.065 -36.305 ;
      RECT -11.165 -36.165 -11.065 -36.065 ;
      RECT -11.165 -35.215 -11.065 -35.115 ;
      RECT -11.165 -31.405 -11.065 -31.305 ;
      RECT -11.165 -30.065 -11.065 -29.965 ;
      RECT -11.165 -26.255 -11.065 -26.155 ;
      RECT -11.165 -25.305 -11.065 -25.205 ;
      RECT -11.165 -25.065 -11.065 -24.965 ;
      RECT -11.165 -23.485 -11.065 -23.385 ;
      RECT -11.165 -23.245 -11.065 -23.145 ;
      RECT -11.165 -22.295 -11.065 -22.195 ;
      RECT -11.165 -18.485 -11.065 -18.385 ;
      RECT -11.165 -17.145 -11.065 -17.045 ;
      RECT -11.165 -13.335 -11.065 -13.235 ;
      RECT -11.165 -12.385 -11.065 -12.285 ;
      RECT -11.165 -12.145 -11.065 -12.045 ;
      RECT -11.165 -10.565 -11.065 -10.465 ;
      RECT -11.165 -10.325 -11.065 -10.225 ;
      RECT -11.165 -9.375 -11.065 -9.275 ;
      RECT -11.165 -5.565 -11.065 -5.465 ;
      RECT -11.165 -4.225 -11.065 -4.125 ;
      RECT -11.165 -0.415 -11.065 -0.315 ;
      RECT -11.165 0.535 -11.065 0.635 ;
      RECT -11.165 0.775 -11.065 0.875 ;
      RECT -11.225 -51.655 -11.125 -51.555 ;
      RECT -11.265 -58.885 -11.165 -58.785 ;
      RECT -11.265 -58.645 -11.165 -58.545 ;
      RECT -11.265 -57.245 -11.165 -57.145 ;
      RECT -11.685 -49.325 -11.585 -49.225 ;
      RECT -11.685 -49.085 -11.585 -48.985 ;
      RECT -11.685 -48.795 -11.585 -48.695 ;
      RECT -11.685 -44.565 -11.585 -44.465 ;
      RECT -11.685 -44.325 -11.585 -44.225 ;
      RECT -11.685 -42.985 -11.585 -42.885 ;
      RECT -11.685 -42.745 -11.585 -42.645 ;
      RECT -11.685 -38.515 -11.585 -38.415 ;
      RECT -11.685 -38.225 -11.585 -38.125 ;
      RECT -11.685 -37.985 -11.585 -37.885 ;
      RECT -11.685 -36.405 -11.585 -36.305 ;
      RECT -11.685 -36.165 -11.585 -36.065 ;
      RECT -11.685 -35.875 -11.585 -35.775 ;
      RECT -11.685 -31.645 -11.585 -31.545 ;
      RECT -11.685 -31.405 -11.585 -31.305 ;
      RECT -11.685 -30.065 -11.585 -29.965 ;
      RECT -11.685 -29.825 -11.585 -29.725 ;
      RECT -11.685 -25.595 -11.585 -25.495 ;
      RECT -11.685 -25.305 -11.585 -25.205 ;
      RECT -11.685 -25.065 -11.585 -24.965 ;
      RECT -11.685 -23.485 -11.585 -23.385 ;
      RECT -11.685 -23.245 -11.585 -23.145 ;
      RECT -11.685 -22.955 -11.585 -22.855 ;
      RECT -11.685 -18.725 -11.585 -18.625 ;
      RECT -11.685 -18.485 -11.585 -18.385 ;
      RECT -11.685 -17.145 -11.585 -17.045 ;
      RECT -11.685 -16.905 -11.585 -16.805 ;
      RECT -11.685 -12.675 -11.585 -12.575 ;
      RECT -11.685 -12.385 -11.585 -12.285 ;
      RECT -11.685 -12.145 -11.585 -12.045 ;
      RECT -11.685 -10.565 -11.585 -10.465 ;
      RECT -11.685 -10.325 -11.585 -10.225 ;
      RECT -11.685 -10.035 -11.585 -9.935 ;
      RECT -11.685 -5.805 -11.585 -5.705 ;
      RECT -11.685 -5.565 -11.585 -5.465 ;
      RECT -11.685 -4.225 -11.585 -4.125 ;
      RECT -11.685 -3.985 -11.585 -3.885 ;
      RECT -11.685 0.245 -11.585 0.345 ;
      RECT -11.685 0.535 -11.585 0.635 ;
      RECT -11.685 0.775 -11.585 0.875 ;
      RECT -11.825 -52.095 -11.725 -51.995 ;
      RECT -11.865 -58.885 -11.765 -58.785 ;
      RECT -11.865 -58.645 -11.765 -58.545 ;
      RECT -11.865 -57.245 -11.765 -57.145 ;
      RECT -12.465 -49.325 -12.365 -49.225 ;
      RECT -12.465 -49.085 -12.365 -48.985 ;
      RECT -12.465 -47.035 -12.365 -46.935 ;
      RECT -12.465 -44.325 -12.365 -44.225 ;
      RECT -12.465 -42.985 -12.365 -42.885 ;
      RECT -12.465 -40.275 -12.365 -40.175 ;
      RECT -12.465 -38.225 -12.365 -38.125 ;
      RECT -12.465 -37.985 -12.365 -37.885 ;
      RECT -12.465 -36.405 -12.365 -36.305 ;
      RECT -12.465 -36.165 -12.365 -36.065 ;
      RECT -12.465 -34.115 -12.365 -34.015 ;
      RECT -12.465 -31.405 -12.365 -31.305 ;
      RECT -12.465 -30.065 -12.365 -29.965 ;
      RECT -12.465 -27.355 -12.365 -27.255 ;
      RECT -12.465 -25.305 -12.365 -25.205 ;
      RECT -12.465 -25.065 -12.365 -24.965 ;
      RECT -12.465 -23.485 -12.365 -23.385 ;
      RECT -12.465 -23.245 -12.365 -23.145 ;
      RECT -12.465 -21.195 -12.365 -21.095 ;
      RECT -12.465 -18.485 -12.365 -18.385 ;
      RECT -12.465 -17.145 -12.365 -17.045 ;
      RECT -12.465 -14.435 -12.365 -14.335 ;
      RECT -12.465 -12.385 -12.365 -12.285 ;
      RECT -12.465 -12.145 -12.365 -12.045 ;
      RECT -12.465 -10.565 -12.365 -10.465 ;
      RECT -12.465 -10.325 -12.365 -10.225 ;
      RECT -12.465 -8.275 -12.365 -8.175 ;
      RECT -12.465 -5.565 -12.365 -5.465 ;
      RECT -12.465 -4.225 -12.365 -4.125 ;
      RECT -12.465 -1.515 -12.365 -1.415 ;
      RECT -12.465 0.535 -12.365 0.635 ;
      RECT -12.465 0.775 -12.365 0.875 ;
      RECT -12.985 -49.325 -12.885 -49.225 ;
      RECT -12.985 -49.085 -12.885 -48.985 ;
      RECT -12.985 -48.795 -12.885 -48.695 ;
      RECT -12.985 -44.565 -12.885 -44.465 ;
      RECT -12.985 -44.325 -12.885 -44.225 ;
      RECT -12.985 -42.985 -12.885 -42.885 ;
      RECT -12.985 -42.745 -12.885 -42.645 ;
      RECT -12.985 -38.515 -12.885 -38.415 ;
      RECT -12.985 -38.225 -12.885 -38.125 ;
      RECT -12.985 -37.985 -12.885 -37.885 ;
      RECT -12.985 -36.405 -12.885 -36.305 ;
      RECT -12.985 -36.165 -12.885 -36.065 ;
      RECT -12.985 -35.875 -12.885 -35.775 ;
      RECT -12.985 -31.645 -12.885 -31.545 ;
      RECT -12.985 -31.405 -12.885 -31.305 ;
      RECT -12.985 -30.065 -12.885 -29.965 ;
      RECT -12.985 -29.825 -12.885 -29.725 ;
      RECT -12.985 -25.595 -12.885 -25.495 ;
      RECT -12.985 -25.305 -12.885 -25.205 ;
      RECT -12.985 -25.065 -12.885 -24.965 ;
      RECT -12.985 -23.485 -12.885 -23.385 ;
      RECT -12.985 -23.245 -12.885 -23.145 ;
      RECT -12.985 -22.955 -12.885 -22.855 ;
      RECT -12.985 -18.725 -12.885 -18.625 ;
      RECT -12.985 -18.485 -12.885 -18.385 ;
      RECT -12.985 -17.145 -12.885 -17.045 ;
      RECT -12.985 -16.905 -12.885 -16.805 ;
      RECT -12.985 -12.675 -12.885 -12.575 ;
      RECT -12.985 -12.385 -12.885 -12.285 ;
      RECT -12.985 -12.145 -12.885 -12.045 ;
      RECT -12.985 -10.565 -12.885 -10.465 ;
      RECT -12.985 -10.325 -12.885 -10.225 ;
      RECT -12.985 -10.035 -12.885 -9.935 ;
      RECT -12.985 -5.805 -12.885 -5.705 ;
      RECT -12.985 -5.565 -12.885 -5.465 ;
      RECT -12.985 -4.225 -12.885 -4.125 ;
      RECT -12.985 -3.985 -12.885 -3.885 ;
      RECT -12.985 0.245 -12.885 0.345 ;
      RECT -12.985 0.535 -12.885 0.635 ;
      RECT -12.985 0.775 -12.885 0.875 ;
      RECT -13.765 -49.325 -13.665 -49.225 ;
      RECT -13.765 -49.085 -13.665 -48.985 ;
      RECT -13.765 -46.815 -13.665 -46.715 ;
      RECT -13.765 -44.325 -13.665 -44.225 ;
      RECT -13.765 -42.985 -13.665 -42.885 ;
      RECT -13.765 -40.495 -13.665 -40.395 ;
      RECT -13.765 -38.225 -13.665 -38.125 ;
      RECT -13.765 -37.985 -13.665 -37.885 ;
      RECT -13.765 -36.405 -13.665 -36.305 ;
      RECT -13.765 -36.165 -13.665 -36.065 ;
      RECT -13.765 -33.895 -13.665 -33.795 ;
      RECT -13.765 -31.405 -13.665 -31.305 ;
      RECT -13.765 -30.065 -13.665 -29.965 ;
      RECT -13.765 -27.575 -13.665 -27.475 ;
      RECT -13.765 -25.305 -13.665 -25.205 ;
      RECT -13.765 -25.065 -13.665 -24.965 ;
      RECT -13.765 -23.485 -13.665 -23.385 ;
      RECT -13.765 -23.245 -13.665 -23.145 ;
      RECT -13.765 -20.975 -13.665 -20.875 ;
      RECT -13.765 -18.485 -13.665 -18.385 ;
      RECT -13.765 -17.145 -13.665 -17.045 ;
      RECT -13.765 -14.655 -13.665 -14.555 ;
      RECT -13.765 -12.385 -13.665 -12.285 ;
      RECT -13.765 -12.145 -13.665 -12.045 ;
      RECT -13.765 -10.565 -13.665 -10.465 ;
      RECT -13.765 -10.325 -13.665 -10.225 ;
      RECT -13.765 -8.055 -13.665 -7.955 ;
      RECT -13.765 -5.565 -13.665 -5.465 ;
      RECT -13.765 -4.225 -13.665 -4.125 ;
      RECT -13.765 -1.735 -13.665 -1.635 ;
      RECT -13.765 0.535 -13.665 0.635 ;
      RECT -13.765 0.775 -13.665 0.875 ;
      RECT -14.285 -49.325 -14.185 -49.225 ;
      RECT -14.285 -49.085 -14.185 -48.985 ;
      RECT -14.285 -48.795 -14.185 -48.695 ;
      RECT -14.285 -44.565 -14.185 -44.465 ;
      RECT -14.285 -44.325 -14.185 -44.225 ;
      RECT -14.285 -42.985 -14.185 -42.885 ;
      RECT -14.285 -42.745 -14.185 -42.645 ;
      RECT -14.285 -38.515 -14.185 -38.415 ;
      RECT -14.285 -38.225 -14.185 -38.125 ;
      RECT -14.285 -37.985 -14.185 -37.885 ;
      RECT -14.285 -36.405 -14.185 -36.305 ;
      RECT -14.285 -36.165 -14.185 -36.065 ;
      RECT -14.285 -35.875 -14.185 -35.775 ;
      RECT -14.285 -31.645 -14.185 -31.545 ;
      RECT -14.285 -31.405 -14.185 -31.305 ;
      RECT -14.285 -30.065 -14.185 -29.965 ;
      RECT -14.285 -29.825 -14.185 -29.725 ;
      RECT -14.285 -25.595 -14.185 -25.495 ;
      RECT -14.285 -25.305 -14.185 -25.205 ;
      RECT -14.285 -25.065 -14.185 -24.965 ;
      RECT -14.285 -23.485 -14.185 -23.385 ;
      RECT -14.285 -23.245 -14.185 -23.145 ;
      RECT -14.285 -22.955 -14.185 -22.855 ;
      RECT -14.285 -18.725 -14.185 -18.625 ;
      RECT -14.285 -18.485 -14.185 -18.385 ;
      RECT -14.285 -17.145 -14.185 -17.045 ;
      RECT -14.285 -16.905 -14.185 -16.805 ;
      RECT -14.285 -12.675 -14.185 -12.575 ;
      RECT -14.285 -12.385 -14.185 -12.285 ;
      RECT -14.285 -12.145 -14.185 -12.045 ;
      RECT -14.285 -10.565 -14.185 -10.465 ;
      RECT -14.285 -10.325 -14.185 -10.225 ;
      RECT -14.285 -10.035 -14.185 -9.935 ;
      RECT -14.285 -5.805 -14.185 -5.705 ;
      RECT -14.285 -5.565 -14.185 -5.465 ;
      RECT -14.285 -4.225 -14.185 -4.125 ;
      RECT -14.285 -3.985 -14.185 -3.885 ;
      RECT -14.285 0.245 -14.185 0.345 ;
      RECT -14.285 0.535 -14.185 0.635 ;
      RECT -14.285 0.775 -14.185 0.875 ;
      RECT -15.065 -49.325 -14.965 -49.225 ;
      RECT -15.065 -49.085 -14.965 -48.985 ;
      RECT -15.065 -47.035 -14.965 -46.935 ;
      RECT -15.065 -44.325 -14.965 -44.225 ;
      RECT -15.065 -42.985 -14.965 -42.885 ;
      RECT -15.065 -40.275 -14.965 -40.175 ;
      RECT -15.065 -38.225 -14.965 -38.125 ;
      RECT -15.065 -37.985 -14.965 -37.885 ;
      RECT -15.065 -36.405 -14.965 -36.305 ;
      RECT -15.065 -36.165 -14.965 -36.065 ;
      RECT -15.065 -34.115 -14.965 -34.015 ;
      RECT -15.065 -31.405 -14.965 -31.305 ;
      RECT -15.065 -30.065 -14.965 -29.965 ;
      RECT -15.065 -27.355 -14.965 -27.255 ;
      RECT -15.065 -25.305 -14.965 -25.205 ;
      RECT -15.065 -25.065 -14.965 -24.965 ;
      RECT -15.065 -23.485 -14.965 -23.385 ;
      RECT -15.065 -23.245 -14.965 -23.145 ;
      RECT -15.065 -21.195 -14.965 -21.095 ;
      RECT -15.065 -18.485 -14.965 -18.385 ;
      RECT -15.065 -17.145 -14.965 -17.045 ;
      RECT -15.065 -14.435 -14.965 -14.335 ;
      RECT -15.065 -12.385 -14.965 -12.285 ;
      RECT -15.065 -12.145 -14.965 -12.045 ;
      RECT -15.065 -10.565 -14.965 -10.465 ;
      RECT -15.065 -10.325 -14.965 -10.225 ;
      RECT -15.065 -8.275 -14.965 -8.175 ;
      RECT -15.065 -5.565 -14.965 -5.465 ;
      RECT -15.065 -4.225 -14.965 -4.125 ;
      RECT -15.065 -1.515 -14.965 -1.415 ;
      RECT -15.065 0.535 -14.965 0.635 ;
      RECT -15.065 0.775 -14.965 0.875 ;
      RECT -15.585 -49.325 -15.485 -49.225 ;
      RECT -15.585 -49.085 -15.485 -48.985 ;
      RECT -15.585 -48.795 -15.485 -48.695 ;
      RECT -15.585 -44.565 -15.485 -44.465 ;
      RECT -15.585 -44.325 -15.485 -44.225 ;
      RECT -15.585 -42.985 -15.485 -42.885 ;
      RECT -15.585 -42.745 -15.485 -42.645 ;
      RECT -15.585 -38.515 -15.485 -38.415 ;
      RECT -15.585 -38.225 -15.485 -38.125 ;
      RECT -15.585 -37.985 -15.485 -37.885 ;
      RECT -15.585 -36.405 -15.485 -36.305 ;
      RECT -15.585 -36.165 -15.485 -36.065 ;
      RECT -15.585 -35.875 -15.485 -35.775 ;
      RECT -15.585 -31.645 -15.485 -31.545 ;
      RECT -15.585 -31.405 -15.485 -31.305 ;
      RECT -15.585 -30.065 -15.485 -29.965 ;
      RECT -15.585 -29.825 -15.485 -29.725 ;
      RECT -15.585 -25.595 -15.485 -25.495 ;
      RECT -15.585 -25.305 -15.485 -25.205 ;
      RECT -15.585 -25.065 -15.485 -24.965 ;
      RECT -15.585 -23.485 -15.485 -23.385 ;
      RECT -15.585 -23.245 -15.485 -23.145 ;
      RECT -15.585 -22.955 -15.485 -22.855 ;
      RECT -15.585 -18.725 -15.485 -18.625 ;
      RECT -15.585 -18.485 -15.485 -18.385 ;
      RECT -15.585 -17.145 -15.485 -17.045 ;
      RECT -15.585 -16.905 -15.485 -16.805 ;
      RECT -15.585 -12.675 -15.485 -12.575 ;
      RECT -15.585 -12.385 -15.485 -12.285 ;
      RECT -15.585 -12.145 -15.485 -12.045 ;
      RECT -15.585 -10.565 -15.485 -10.465 ;
      RECT -15.585 -10.325 -15.485 -10.225 ;
      RECT -15.585 -10.035 -15.485 -9.935 ;
      RECT -15.585 -5.805 -15.485 -5.705 ;
      RECT -15.585 -5.565 -15.485 -5.465 ;
      RECT -15.585 -4.225 -15.485 -4.125 ;
      RECT -15.585 -3.985 -15.485 -3.885 ;
      RECT -15.585 0.245 -15.485 0.345 ;
      RECT -15.585 0.535 -15.485 0.635 ;
      RECT -15.585 0.775 -15.485 0.875 ;
      RECT -16.365 -49.325 -16.265 -49.225 ;
      RECT -16.365 -49.085 -16.265 -48.985 ;
      RECT -16.365 -46.375 -16.265 -46.275 ;
      RECT -16.365 -44.325 -16.265 -44.225 ;
      RECT -16.365 -42.985 -16.265 -42.885 ;
      RECT -16.365 -40.935 -16.265 -40.835 ;
      RECT -16.365 -38.225 -16.265 -38.125 ;
      RECT -16.365 -37.985 -16.265 -37.885 ;
      RECT -16.365 -36.405 -16.265 -36.305 ;
      RECT -16.365 -36.165 -16.265 -36.065 ;
      RECT -16.365 -33.455 -16.265 -33.355 ;
      RECT -16.365 -31.405 -16.265 -31.305 ;
      RECT -16.365 -30.065 -16.265 -29.965 ;
      RECT -16.365 -28.015 -16.265 -27.915 ;
      RECT -16.365 -25.305 -16.265 -25.205 ;
      RECT -16.365 -25.065 -16.265 -24.965 ;
      RECT -16.365 -23.485 -16.265 -23.385 ;
      RECT -16.365 -23.245 -16.265 -23.145 ;
      RECT -16.365 -20.535 -16.265 -20.435 ;
      RECT -16.365 -18.485 -16.265 -18.385 ;
      RECT -16.365 -17.145 -16.265 -17.045 ;
      RECT -16.365 -15.095 -16.265 -14.995 ;
      RECT -16.365 -12.385 -16.265 -12.285 ;
      RECT -16.365 -12.145 -16.265 -12.045 ;
      RECT -16.365 -10.565 -16.265 -10.465 ;
      RECT -16.365 -10.325 -16.265 -10.225 ;
      RECT -16.365 -7.615 -16.265 -7.515 ;
      RECT -16.365 -5.565 -16.265 -5.465 ;
      RECT -16.365 -4.225 -16.265 -4.125 ;
      RECT -16.365 -2.175 -16.265 -2.075 ;
      RECT -16.365 0.535 -16.265 0.635 ;
      RECT -16.365 0.775 -16.265 0.875 ;
      RECT -16.885 -49.325 -16.785 -49.225 ;
      RECT -16.885 -49.085 -16.785 -48.985 ;
      RECT -16.885 -48.795 -16.785 -48.695 ;
      RECT -16.885 -44.565 -16.785 -44.465 ;
      RECT -16.885 -44.325 -16.785 -44.225 ;
      RECT -16.885 -42.985 -16.785 -42.885 ;
      RECT -16.885 -42.745 -16.785 -42.645 ;
      RECT -16.885 -38.515 -16.785 -38.415 ;
      RECT -16.885 -38.225 -16.785 -38.125 ;
      RECT -16.885 -37.985 -16.785 -37.885 ;
      RECT -16.885 -36.405 -16.785 -36.305 ;
      RECT -16.885 -36.165 -16.785 -36.065 ;
      RECT -16.885 -35.875 -16.785 -35.775 ;
      RECT -16.885 -31.645 -16.785 -31.545 ;
      RECT -16.885 -31.405 -16.785 -31.305 ;
      RECT -16.885 -30.065 -16.785 -29.965 ;
      RECT -16.885 -29.825 -16.785 -29.725 ;
      RECT -16.885 -25.595 -16.785 -25.495 ;
      RECT -16.885 -25.305 -16.785 -25.205 ;
      RECT -16.885 -25.065 -16.785 -24.965 ;
      RECT -16.885 -23.485 -16.785 -23.385 ;
      RECT -16.885 -23.245 -16.785 -23.145 ;
      RECT -16.885 -22.955 -16.785 -22.855 ;
      RECT -16.885 -18.725 -16.785 -18.625 ;
      RECT -16.885 -18.485 -16.785 -18.385 ;
      RECT -16.885 -17.145 -16.785 -17.045 ;
      RECT -16.885 -16.905 -16.785 -16.805 ;
      RECT -16.885 -12.675 -16.785 -12.575 ;
      RECT -16.885 -12.385 -16.785 -12.285 ;
      RECT -16.885 -12.145 -16.785 -12.045 ;
      RECT -16.885 -10.565 -16.785 -10.465 ;
      RECT -16.885 -10.325 -16.785 -10.225 ;
      RECT -16.885 -10.035 -16.785 -9.935 ;
      RECT -16.885 -5.805 -16.785 -5.705 ;
      RECT -16.885 -5.565 -16.785 -5.465 ;
      RECT -16.885 -4.225 -16.785 -4.125 ;
      RECT -16.885 -3.985 -16.785 -3.885 ;
      RECT -16.885 0.245 -16.785 0.345 ;
      RECT -16.885 0.535 -16.785 0.635 ;
      RECT -16.885 0.775 -16.785 0.875 ;
      RECT -17.665 -49.325 -17.565 -49.225 ;
      RECT -17.665 -49.085 -17.565 -48.985 ;
      RECT -17.665 -47.035 -17.565 -46.935 ;
      RECT -17.665 -44.325 -17.565 -44.225 ;
      RECT -17.665 -42.985 -17.565 -42.885 ;
      RECT -17.665 -40.275 -17.565 -40.175 ;
      RECT -17.665 -38.225 -17.565 -38.125 ;
      RECT -17.665 -37.985 -17.565 -37.885 ;
      RECT -17.665 -36.405 -17.565 -36.305 ;
      RECT -17.665 -36.165 -17.565 -36.065 ;
      RECT -17.665 -34.115 -17.565 -34.015 ;
      RECT -17.665 -31.405 -17.565 -31.305 ;
      RECT -17.665 -30.065 -17.565 -29.965 ;
      RECT -17.665 -27.355 -17.565 -27.255 ;
      RECT -17.665 -25.305 -17.565 -25.205 ;
      RECT -17.665 -25.065 -17.565 -24.965 ;
      RECT -17.665 -23.485 -17.565 -23.385 ;
      RECT -17.665 -23.245 -17.565 -23.145 ;
      RECT -17.665 -21.195 -17.565 -21.095 ;
      RECT -17.665 -18.485 -17.565 -18.385 ;
      RECT -17.665 -17.145 -17.565 -17.045 ;
      RECT -17.665 -14.435 -17.565 -14.335 ;
      RECT -17.665 -12.385 -17.565 -12.285 ;
      RECT -17.665 -12.145 -17.565 -12.045 ;
      RECT -17.665 -10.565 -17.565 -10.465 ;
      RECT -17.665 -10.325 -17.565 -10.225 ;
      RECT -17.665 -8.275 -17.565 -8.175 ;
      RECT -17.665 -5.565 -17.565 -5.465 ;
      RECT -17.665 -4.225 -17.565 -4.125 ;
      RECT -17.665 -1.515 -17.565 -1.415 ;
      RECT -17.665 0.535 -17.565 0.635 ;
      RECT -17.665 0.775 -17.565 0.875 ;
      RECT -18.185 -49.325 -18.085 -49.225 ;
      RECT -18.185 -49.085 -18.085 -48.985 ;
      RECT -18.185 -48.795 -18.085 -48.695 ;
      RECT -18.185 -44.565 -18.085 -44.465 ;
      RECT -18.185 -44.325 -18.085 -44.225 ;
      RECT -18.185 -42.985 -18.085 -42.885 ;
      RECT -18.185 -42.745 -18.085 -42.645 ;
      RECT -18.185 -38.515 -18.085 -38.415 ;
      RECT -18.185 -38.225 -18.085 -38.125 ;
      RECT -18.185 -37.985 -18.085 -37.885 ;
      RECT -18.185 -36.405 -18.085 -36.305 ;
      RECT -18.185 -36.165 -18.085 -36.065 ;
      RECT -18.185 -35.875 -18.085 -35.775 ;
      RECT -18.185 -31.645 -18.085 -31.545 ;
      RECT -18.185 -31.405 -18.085 -31.305 ;
      RECT -18.185 -30.065 -18.085 -29.965 ;
      RECT -18.185 -29.825 -18.085 -29.725 ;
      RECT -18.185 -25.595 -18.085 -25.495 ;
      RECT -18.185 -25.305 -18.085 -25.205 ;
      RECT -18.185 -25.065 -18.085 -24.965 ;
      RECT -18.185 -23.485 -18.085 -23.385 ;
      RECT -18.185 -23.245 -18.085 -23.145 ;
      RECT -18.185 -22.955 -18.085 -22.855 ;
      RECT -18.185 -18.725 -18.085 -18.625 ;
      RECT -18.185 -18.485 -18.085 -18.385 ;
      RECT -18.185 -17.145 -18.085 -17.045 ;
      RECT -18.185 -16.905 -18.085 -16.805 ;
      RECT -18.185 -12.675 -18.085 -12.575 ;
      RECT -18.185 -12.385 -18.085 -12.285 ;
      RECT -18.185 -12.145 -18.085 -12.045 ;
      RECT -18.185 -10.565 -18.085 -10.465 ;
      RECT -18.185 -10.325 -18.085 -10.225 ;
      RECT -18.185 -10.035 -18.085 -9.935 ;
      RECT -18.185 -5.805 -18.085 -5.705 ;
      RECT -18.185 -5.565 -18.085 -5.465 ;
      RECT -18.185 -4.225 -18.085 -4.125 ;
      RECT -18.185 -3.985 -18.085 -3.885 ;
      RECT -18.185 0.245 -18.085 0.345 ;
      RECT -18.185 0.535 -18.085 0.635 ;
      RECT -18.185 0.775 -18.085 0.875 ;
      RECT -18.965 -49.325 -18.865 -49.225 ;
      RECT -18.965 -49.085 -18.865 -48.985 ;
      RECT -18.965 -46.815 -18.865 -46.715 ;
      RECT -18.965 -44.325 -18.865 -44.225 ;
      RECT -18.965 -42.985 -18.865 -42.885 ;
      RECT -18.965 -40.495 -18.865 -40.395 ;
      RECT -18.965 -38.225 -18.865 -38.125 ;
      RECT -18.965 -37.985 -18.865 -37.885 ;
      RECT -18.965 -36.405 -18.865 -36.305 ;
      RECT -18.965 -36.165 -18.865 -36.065 ;
      RECT -18.965 -33.895 -18.865 -33.795 ;
      RECT -18.965 -31.405 -18.865 -31.305 ;
      RECT -18.965 -30.065 -18.865 -29.965 ;
      RECT -18.965 -27.575 -18.865 -27.475 ;
      RECT -18.965 -25.305 -18.865 -25.205 ;
      RECT -18.965 -25.065 -18.865 -24.965 ;
      RECT -18.965 -23.485 -18.865 -23.385 ;
      RECT -18.965 -23.245 -18.865 -23.145 ;
      RECT -18.965 -20.975 -18.865 -20.875 ;
      RECT -18.965 -18.485 -18.865 -18.385 ;
      RECT -18.965 -17.145 -18.865 -17.045 ;
      RECT -18.965 -14.655 -18.865 -14.555 ;
      RECT -18.965 -12.385 -18.865 -12.285 ;
      RECT -18.965 -12.145 -18.865 -12.045 ;
      RECT -18.965 -10.565 -18.865 -10.465 ;
      RECT -18.965 -10.325 -18.865 -10.225 ;
      RECT -18.965 -8.055 -18.865 -7.955 ;
      RECT -18.965 -5.565 -18.865 -5.465 ;
      RECT -18.965 -4.225 -18.865 -4.125 ;
      RECT -18.965 -1.735 -18.865 -1.635 ;
      RECT -18.965 0.535 -18.865 0.635 ;
      RECT -18.965 0.775 -18.865 0.875 ;
      RECT -19.485 -49.325 -19.385 -49.225 ;
      RECT -19.485 -49.085 -19.385 -48.985 ;
      RECT -19.485 -48.795 -19.385 -48.695 ;
      RECT -19.485 -44.565 -19.385 -44.465 ;
      RECT -19.485 -44.325 -19.385 -44.225 ;
      RECT -19.485 -42.985 -19.385 -42.885 ;
      RECT -19.485 -42.745 -19.385 -42.645 ;
      RECT -19.485 -38.515 -19.385 -38.415 ;
      RECT -19.485 -38.225 -19.385 -38.125 ;
      RECT -19.485 -37.985 -19.385 -37.885 ;
      RECT -19.485 -36.405 -19.385 -36.305 ;
      RECT -19.485 -36.165 -19.385 -36.065 ;
      RECT -19.485 -35.875 -19.385 -35.775 ;
      RECT -19.485 -31.645 -19.385 -31.545 ;
      RECT -19.485 -31.405 -19.385 -31.305 ;
      RECT -19.485 -30.065 -19.385 -29.965 ;
      RECT -19.485 -29.825 -19.385 -29.725 ;
      RECT -19.485 -25.595 -19.385 -25.495 ;
      RECT -19.485 -25.305 -19.385 -25.205 ;
      RECT -19.485 -25.065 -19.385 -24.965 ;
      RECT -19.485 -23.485 -19.385 -23.385 ;
      RECT -19.485 -23.245 -19.385 -23.145 ;
      RECT -19.485 -22.955 -19.385 -22.855 ;
      RECT -19.485 -18.725 -19.385 -18.625 ;
      RECT -19.485 -18.485 -19.385 -18.385 ;
      RECT -19.485 -17.145 -19.385 -17.045 ;
      RECT -19.485 -16.905 -19.385 -16.805 ;
      RECT -19.485 -12.675 -19.385 -12.575 ;
      RECT -19.485 -12.385 -19.385 -12.285 ;
      RECT -19.485 -12.145 -19.385 -12.045 ;
      RECT -19.485 -10.565 -19.385 -10.465 ;
      RECT -19.485 -10.325 -19.385 -10.225 ;
      RECT -19.485 -10.035 -19.385 -9.935 ;
      RECT -19.485 -5.805 -19.385 -5.705 ;
      RECT -19.485 -5.565 -19.385 -5.465 ;
      RECT -19.485 -4.225 -19.385 -4.125 ;
      RECT -19.485 -3.985 -19.385 -3.885 ;
      RECT -19.485 0.245 -19.385 0.345 ;
      RECT -19.485 0.535 -19.385 0.635 ;
      RECT -19.485 0.775 -19.385 0.875 ;
      RECT -20.265 -49.325 -20.165 -49.225 ;
      RECT -20.265 -49.085 -20.165 -48.985 ;
      RECT -20.265 -47.035 -20.165 -46.935 ;
      RECT -20.265 -44.325 -20.165 -44.225 ;
      RECT -20.265 -42.985 -20.165 -42.885 ;
      RECT -20.265 -40.275 -20.165 -40.175 ;
      RECT -20.265 -38.225 -20.165 -38.125 ;
      RECT -20.265 -37.985 -20.165 -37.885 ;
      RECT -20.265 -36.405 -20.165 -36.305 ;
      RECT -20.265 -36.165 -20.165 -36.065 ;
      RECT -20.265 -34.115 -20.165 -34.015 ;
      RECT -20.265 -31.405 -20.165 -31.305 ;
      RECT -20.265 -30.065 -20.165 -29.965 ;
      RECT -20.265 -27.355 -20.165 -27.255 ;
      RECT -20.265 -25.305 -20.165 -25.205 ;
      RECT -20.265 -25.065 -20.165 -24.965 ;
      RECT -20.265 -23.485 -20.165 -23.385 ;
      RECT -20.265 -23.245 -20.165 -23.145 ;
      RECT -20.265 -21.195 -20.165 -21.095 ;
      RECT -20.265 -18.485 -20.165 -18.385 ;
      RECT -20.265 -17.145 -20.165 -17.045 ;
      RECT -20.265 -14.435 -20.165 -14.335 ;
      RECT -20.265 -12.385 -20.165 -12.285 ;
      RECT -20.265 -12.145 -20.165 -12.045 ;
      RECT -20.265 -10.565 -20.165 -10.465 ;
      RECT -20.265 -10.325 -20.165 -10.225 ;
      RECT -20.265 -8.275 -20.165 -8.175 ;
      RECT -20.265 -5.565 -20.165 -5.465 ;
      RECT -20.265 -4.225 -20.165 -4.125 ;
      RECT -20.265 -1.515 -20.165 -1.415 ;
      RECT -20.265 0.535 -20.165 0.635 ;
      RECT -20.265 0.775 -20.165 0.875 ;
      RECT -20.785 -49.325 -20.685 -49.225 ;
      RECT -20.785 -49.085 -20.685 -48.985 ;
      RECT -20.785 -48.795 -20.685 -48.695 ;
      RECT -20.785 -44.565 -20.685 -44.465 ;
      RECT -20.785 -44.325 -20.685 -44.225 ;
      RECT -20.785 -42.985 -20.685 -42.885 ;
      RECT -20.785 -42.745 -20.685 -42.645 ;
      RECT -20.785 -38.515 -20.685 -38.415 ;
      RECT -20.785 -38.225 -20.685 -38.125 ;
      RECT -20.785 -37.985 -20.685 -37.885 ;
      RECT -20.785 -36.405 -20.685 -36.305 ;
      RECT -20.785 -36.165 -20.685 -36.065 ;
      RECT -20.785 -35.875 -20.685 -35.775 ;
      RECT -20.785 -31.645 -20.685 -31.545 ;
      RECT -20.785 -31.405 -20.685 -31.305 ;
      RECT -20.785 -30.065 -20.685 -29.965 ;
      RECT -20.785 -29.825 -20.685 -29.725 ;
      RECT -20.785 -25.595 -20.685 -25.495 ;
      RECT -20.785 -25.305 -20.685 -25.205 ;
      RECT -20.785 -25.065 -20.685 -24.965 ;
      RECT -20.785 -23.485 -20.685 -23.385 ;
      RECT -20.785 -23.245 -20.685 -23.145 ;
      RECT -20.785 -22.955 -20.685 -22.855 ;
      RECT -20.785 -18.725 -20.685 -18.625 ;
      RECT -20.785 -18.485 -20.685 -18.385 ;
      RECT -20.785 -17.145 -20.685 -17.045 ;
      RECT -20.785 -16.905 -20.685 -16.805 ;
      RECT -20.785 -12.675 -20.685 -12.575 ;
      RECT -20.785 -12.385 -20.685 -12.285 ;
      RECT -20.785 -12.145 -20.685 -12.045 ;
      RECT -20.785 -10.565 -20.685 -10.465 ;
      RECT -20.785 -10.325 -20.685 -10.225 ;
      RECT -20.785 -10.035 -20.685 -9.935 ;
      RECT -20.785 -5.805 -20.685 -5.705 ;
      RECT -20.785 -5.565 -20.685 -5.465 ;
      RECT -20.785 -4.225 -20.685 -4.125 ;
      RECT -20.785 -3.985 -20.685 -3.885 ;
      RECT -20.785 0.245 -20.685 0.345 ;
      RECT -20.785 0.535 -20.685 0.635 ;
      RECT -20.785 0.775 -20.685 0.875 ;
      RECT -21.565 -49.325 -21.465 -49.225 ;
      RECT -21.565 -49.085 -21.465 -48.985 ;
      RECT -21.565 -46.595 -21.465 -46.495 ;
      RECT -21.565 -44.325 -21.465 -44.225 ;
      RECT -21.565 -42.985 -21.465 -42.885 ;
      RECT -21.565 -40.715 -21.465 -40.615 ;
      RECT -21.565 -38.225 -21.465 -38.125 ;
      RECT -21.565 -37.985 -21.465 -37.885 ;
      RECT -21.565 -36.405 -21.465 -36.305 ;
      RECT -21.565 -36.165 -21.465 -36.065 ;
      RECT -21.565 -33.675 -21.465 -33.575 ;
      RECT -21.565 -31.405 -21.465 -31.305 ;
      RECT -21.565 -30.065 -21.465 -29.965 ;
      RECT -21.565 -27.795 -21.465 -27.695 ;
      RECT -21.565 -25.305 -21.465 -25.205 ;
      RECT -21.565 -25.065 -21.465 -24.965 ;
      RECT -21.565 -23.485 -21.465 -23.385 ;
      RECT -21.565 -23.245 -21.465 -23.145 ;
      RECT -21.565 -20.755 -21.465 -20.655 ;
      RECT -21.565 -18.485 -21.465 -18.385 ;
      RECT -21.565 -17.145 -21.465 -17.045 ;
      RECT -21.565 -14.875 -21.465 -14.775 ;
      RECT -21.565 -12.385 -21.465 -12.285 ;
      RECT -21.565 -12.145 -21.465 -12.045 ;
      RECT -21.565 -10.565 -21.465 -10.465 ;
      RECT -21.565 -10.325 -21.465 -10.225 ;
      RECT -21.565 -7.835 -21.465 -7.735 ;
      RECT -21.565 -5.565 -21.465 -5.465 ;
      RECT -21.565 -4.225 -21.465 -4.125 ;
      RECT -21.565 -1.955 -21.465 -1.855 ;
      RECT -21.565 0.535 -21.465 0.635 ;
      RECT -21.565 0.775 -21.465 0.875 ;
      RECT -22.085 -49.325 -21.985 -49.225 ;
      RECT -22.085 -49.085 -21.985 -48.985 ;
      RECT -22.085 -48.795 -21.985 -48.695 ;
      RECT -22.085 -44.565 -21.985 -44.465 ;
      RECT -22.085 -44.325 -21.985 -44.225 ;
      RECT -22.085 -42.985 -21.985 -42.885 ;
      RECT -22.085 -42.745 -21.985 -42.645 ;
      RECT -22.085 -38.515 -21.985 -38.415 ;
      RECT -22.085 -38.225 -21.985 -38.125 ;
      RECT -22.085 -37.985 -21.985 -37.885 ;
      RECT -22.085 -36.405 -21.985 -36.305 ;
      RECT -22.085 -36.165 -21.985 -36.065 ;
      RECT -22.085 -35.875 -21.985 -35.775 ;
      RECT -22.085 -31.645 -21.985 -31.545 ;
      RECT -22.085 -31.405 -21.985 -31.305 ;
      RECT -22.085 -30.065 -21.985 -29.965 ;
      RECT -22.085 -29.825 -21.985 -29.725 ;
      RECT -22.085 -25.595 -21.985 -25.495 ;
      RECT -22.085 -25.305 -21.985 -25.205 ;
      RECT -22.085 -25.065 -21.985 -24.965 ;
      RECT -22.085 -23.485 -21.985 -23.385 ;
      RECT -22.085 -23.245 -21.985 -23.145 ;
      RECT -22.085 -22.955 -21.985 -22.855 ;
      RECT -22.085 -18.725 -21.985 -18.625 ;
      RECT -22.085 -18.485 -21.985 -18.385 ;
      RECT -22.085 -17.145 -21.985 -17.045 ;
      RECT -22.085 -16.905 -21.985 -16.805 ;
      RECT -22.085 -12.675 -21.985 -12.575 ;
      RECT -22.085 -12.385 -21.985 -12.285 ;
      RECT -22.085 -12.145 -21.985 -12.045 ;
      RECT -22.085 -10.565 -21.985 -10.465 ;
      RECT -22.085 -10.325 -21.985 -10.225 ;
      RECT -22.085 -10.035 -21.985 -9.935 ;
      RECT -22.085 -5.805 -21.985 -5.705 ;
      RECT -22.085 -5.565 -21.985 -5.465 ;
      RECT -22.085 -4.225 -21.985 -4.125 ;
      RECT -22.085 -3.985 -21.985 -3.885 ;
      RECT -22.085 0.245 -21.985 0.345 ;
      RECT -22.085 0.535 -21.985 0.635 ;
      RECT -22.085 0.775 -21.985 0.875 ;
      RECT -22.865 -49.325 -22.765 -49.225 ;
      RECT -22.865 -49.085 -22.765 -48.985 ;
      RECT -22.865 -47.035 -22.765 -46.935 ;
      RECT -22.865 -44.325 -22.765 -44.225 ;
      RECT -22.865 -42.985 -22.765 -42.885 ;
      RECT -22.865 -40.275 -22.765 -40.175 ;
      RECT -22.865 -38.225 -22.765 -38.125 ;
      RECT -22.865 -37.985 -22.765 -37.885 ;
      RECT -22.865 -36.405 -22.765 -36.305 ;
      RECT -22.865 -36.165 -22.765 -36.065 ;
      RECT -22.865 -34.115 -22.765 -34.015 ;
      RECT -22.865 -31.405 -22.765 -31.305 ;
      RECT -22.865 -30.065 -22.765 -29.965 ;
      RECT -22.865 -27.355 -22.765 -27.255 ;
      RECT -22.865 -25.305 -22.765 -25.205 ;
      RECT -22.865 -25.065 -22.765 -24.965 ;
      RECT -22.865 -23.485 -22.765 -23.385 ;
      RECT -22.865 -23.245 -22.765 -23.145 ;
      RECT -22.865 -21.195 -22.765 -21.095 ;
      RECT -22.865 -18.485 -22.765 -18.385 ;
      RECT -22.865 -17.145 -22.765 -17.045 ;
      RECT -22.865 -14.435 -22.765 -14.335 ;
      RECT -22.865 -12.385 -22.765 -12.285 ;
      RECT -22.865 -12.145 -22.765 -12.045 ;
      RECT -22.865 -10.565 -22.765 -10.465 ;
      RECT -22.865 -10.325 -22.765 -10.225 ;
      RECT -22.865 -8.275 -22.765 -8.175 ;
      RECT -22.865 -5.565 -22.765 -5.465 ;
      RECT -22.865 -4.225 -22.765 -4.125 ;
      RECT -22.865 -1.515 -22.765 -1.415 ;
      RECT -22.865 0.535 -22.765 0.635 ;
      RECT -22.865 0.775 -22.765 0.875 ;
      RECT -23.385 -49.325 -23.285 -49.225 ;
      RECT -23.385 -49.085 -23.285 -48.985 ;
      RECT -23.385 -48.795 -23.285 -48.695 ;
      RECT -23.385 -44.565 -23.285 -44.465 ;
      RECT -23.385 -44.325 -23.285 -44.225 ;
      RECT -23.385 -42.985 -23.285 -42.885 ;
      RECT -23.385 -42.745 -23.285 -42.645 ;
      RECT -23.385 -38.515 -23.285 -38.415 ;
      RECT -23.385 -38.225 -23.285 -38.125 ;
      RECT -23.385 -37.985 -23.285 -37.885 ;
      RECT -23.385 -36.405 -23.285 -36.305 ;
      RECT -23.385 -36.165 -23.285 -36.065 ;
      RECT -23.385 -35.875 -23.285 -35.775 ;
      RECT -23.385 -31.645 -23.285 -31.545 ;
      RECT -23.385 -31.405 -23.285 -31.305 ;
      RECT -23.385 -30.065 -23.285 -29.965 ;
      RECT -23.385 -29.825 -23.285 -29.725 ;
      RECT -23.385 -25.595 -23.285 -25.495 ;
      RECT -23.385 -25.305 -23.285 -25.205 ;
      RECT -23.385 -25.065 -23.285 -24.965 ;
      RECT -23.385 -23.485 -23.285 -23.385 ;
      RECT -23.385 -23.245 -23.285 -23.145 ;
      RECT -23.385 -22.955 -23.285 -22.855 ;
      RECT -23.385 -18.725 -23.285 -18.625 ;
      RECT -23.385 -18.485 -23.285 -18.385 ;
      RECT -23.385 -17.145 -23.285 -17.045 ;
      RECT -23.385 -16.905 -23.285 -16.805 ;
      RECT -23.385 -12.675 -23.285 -12.575 ;
      RECT -23.385 -12.385 -23.285 -12.285 ;
      RECT -23.385 -12.145 -23.285 -12.045 ;
      RECT -23.385 -10.565 -23.285 -10.465 ;
      RECT -23.385 -10.325 -23.285 -10.225 ;
      RECT -23.385 -10.035 -23.285 -9.935 ;
      RECT -23.385 -5.805 -23.285 -5.705 ;
      RECT -23.385 -5.565 -23.285 -5.465 ;
      RECT -23.385 -4.225 -23.285 -4.125 ;
      RECT -23.385 -3.985 -23.285 -3.885 ;
      RECT -23.385 0.245 -23.285 0.345 ;
      RECT -23.385 0.535 -23.285 0.635 ;
      RECT -23.385 0.775 -23.285 0.875 ;
      RECT -24.165 -49.325 -24.065 -49.225 ;
      RECT -24.165 -49.085 -24.065 -48.985 ;
      RECT -24.165 -46.815 -24.065 -46.715 ;
      RECT -24.165 -44.325 -24.065 -44.225 ;
      RECT -24.165 -42.985 -24.065 -42.885 ;
      RECT -24.165 -40.495 -24.065 -40.395 ;
      RECT -24.165 -38.225 -24.065 -38.125 ;
      RECT -24.165 -37.985 -24.065 -37.885 ;
      RECT -24.165 -36.405 -24.065 -36.305 ;
      RECT -24.165 -36.165 -24.065 -36.065 ;
      RECT -24.165 -33.895 -24.065 -33.795 ;
      RECT -24.165 -31.405 -24.065 -31.305 ;
      RECT -24.165 -30.065 -24.065 -29.965 ;
      RECT -24.165 -27.575 -24.065 -27.475 ;
      RECT -24.165 -25.305 -24.065 -25.205 ;
      RECT -24.165 -25.065 -24.065 -24.965 ;
      RECT -24.165 -23.485 -24.065 -23.385 ;
      RECT -24.165 -23.245 -24.065 -23.145 ;
      RECT -24.165 -20.975 -24.065 -20.875 ;
      RECT -24.165 -18.485 -24.065 -18.385 ;
      RECT -24.165 -17.145 -24.065 -17.045 ;
      RECT -24.165 -14.655 -24.065 -14.555 ;
      RECT -24.165 -12.385 -24.065 -12.285 ;
      RECT -24.165 -12.145 -24.065 -12.045 ;
      RECT -24.165 -10.565 -24.065 -10.465 ;
      RECT -24.165 -10.325 -24.065 -10.225 ;
      RECT -24.165 -8.055 -24.065 -7.955 ;
      RECT -24.165 -5.565 -24.065 -5.465 ;
      RECT -24.165 -4.225 -24.065 -4.125 ;
      RECT -24.165 -1.735 -24.065 -1.635 ;
      RECT -24.165 0.535 -24.065 0.635 ;
      RECT -24.165 0.775 -24.065 0.875 ;
      RECT -24.685 -49.325 -24.585 -49.225 ;
      RECT -24.685 -49.085 -24.585 -48.985 ;
      RECT -24.685 -48.795 -24.585 -48.695 ;
      RECT -24.685 -44.565 -24.585 -44.465 ;
      RECT -24.685 -44.325 -24.585 -44.225 ;
      RECT -24.685 -42.985 -24.585 -42.885 ;
      RECT -24.685 -42.745 -24.585 -42.645 ;
      RECT -24.685 -38.515 -24.585 -38.415 ;
      RECT -24.685 -38.225 -24.585 -38.125 ;
      RECT -24.685 -37.985 -24.585 -37.885 ;
      RECT -24.685 -36.405 -24.585 -36.305 ;
      RECT -24.685 -36.165 -24.585 -36.065 ;
      RECT -24.685 -35.875 -24.585 -35.775 ;
      RECT -24.685 -31.645 -24.585 -31.545 ;
      RECT -24.685 -31.405 -24.585 -31.305 ;
      RECT -24.685 -30.065 -24.585 -29.965 ;
      RECT -24.685 -29.825 -24.585 -29.725 ;
      RECT -24.685 -25.595 -24.585 -25.495 ;
      RECT -24.685 -25.305 -24.585 -25.205 ;
      RECT -24.685 -25.065 -24.585 -24.965 ;
      RECT -24.685 -23.485 -24.585 -23.385 ;
      RECT -24.685 -23.245 -24.585 -23.145 ;
      RECT -24.685 -22.955 -24.585 -22.855 ;
      RECT -24.685 -18.725 -24.585 -18.625 ;
      RECT -24.685 -18.485 -24.585 -18.385 ;
      RECT -24.685 -17.145 -24.585 -17.045 ;
      RECT -24.685 -16.905 -24.585 -16.805 ;
      RECT -24.685 -12.675 -24.585 -12.575 ;
      RECT -24.685 -12.385 -24.585 -12.285 ;
      RECT -24.685 -12.145 -24.585 -12.045 ;
      RECT -24.685 -10.565 -24.585 -10.465 ;
      RECT -24.685 -10.325 -24.585 -10.225 ;
      RECT -24.685 -10.035 -24.585 -9.935 ;
      RECT -24.685 -5.805 -24.585 -5.705 ;
      RECT -24.685 -5.565 -24.585 -5.465 ;
      RECT -24.685 -4.225 -24.585 -4.125 ;
      RECT -24.685 -3.985 -24.585 -3.885 ;
      RECT -24.685 0.245 -24.585 0.345 ;
      RECT -24.685 0.535 -24.585 0.635 ;
      RECT -24.685 0.775 -24.585 0.875 ;
      RECT -25.465 -49.325 -25.365 -49.225 ;
      RECT -25.465 -49.085 -25.365 -48.985 ;
      RECT -25.465 -47.035 -25.365 -46.935 ;
      RECT -25.465 -44.325 -25.365 -44.225 ;
      RECT -25.465 -42.985 -25.365 -42.885 ;
      RECT -25.465 -40.275 -25.365 -40.175 ;
      RECT -25.465 -38.225 -25.365 -38.125 ;
      RECT -25.465 -37.985 -25.365 -37.885 ;
      RECT -25.465 -36.405 -25.365 -36.305 ;
      RECT -25.465 -36.165 -25.365 -36.065 ;
      RECT -25.465 -34.115 -25.365 -34.015 ;
      RECT -25.465 -31.405 -25.365 -31.305 ;
      RECT -25.465 -30.065 -25.365 -29.965 ;
      RECT -25.465 -27.355 -25.365 -27.255 ;
      RECT -25.465 -25.305 -25.365 -25.205 ;
      RECT -25.465 -25.065 -25.365 -24.965 ;
      RECT -25.465 -23.485 -25.365 -23.385 ;
      RECT -25.465 -23.245 -25.365 -23.145 ;
      RECT -25.465 -21.195 -25.365 -21.095 ;
      RECT -25.465 -18.485 -25.365 -18.385 ;
      RECT -25.465 -17.145 -25.365 -17.045 ;
      RECT -25.465 -14.435 -25.365 -14.335 ;
      RECT -25.465 -12.385 -25.365 -12.285 ;
      RECT -25.465 -12.145 -25.365 -12.045 ;
      RECT -25.465 -10.565 -25.365 -10.465 ;
      RECT -25.465 -10.325 -25.365 -10.225 ;
      RECT -25.465 -8.275 -25.365 -8.175 ;
      RECT -25.465 -5.565 -25.365 -5.465 ;
      RECT -25.465 -4.225 -25.365 -4.125 ;
      RECT -25.465 -1.515 -25.365 -1.415 ;
      RECT -25.465 0.535 -25.365 0.635 ;
      RECT -25.465 0.775 -25.365 0.875 ;
      RECT -25.985 -49.325 -25.885 -49.225 ;
      RECT -25.985 -49.085 -25.885 -48.985 ;
      RECT -25.985 -48.795 -25.885 -48.695 ;
      RECT -25.985 -44.565 -25.885 -44.465 ;
      RECT -25.985 -44.325 -25.885 -44.225 ;
      RECT -25.985 -42.985 -25.885 -42.885 ;
      RECT -25.985 -42.745 -25.885 -42.645 ;
      RECT -25.985 -38.515 -25.885 -38.415 ;
      RECT -25.985 -38.225 -25.885 -38.125 ;
      RECT -25.985 -37.985 -25.885 -37.885 ;
      RECT -25.985 -36.405 -25.885 -36.305 ;
      RECT -25.985 -36.165 -25.885 -36.065 ;
      RECT -25.985 -35.875 -25.885 -35.775 ;
      RECT -25.985 -31.645 -25.885 -31.545 ;
      RECT -25.985 -31.405 -25.885 -31.305 ;
      RECT -25.985 -30.065 -25.885 -29.965 ;
      RECT -25.985 -29.825 -25.885 -29.725 ;
      RECT -25.985 -25.595 -25.885 -25.495 ;
      RECT -25.985 -25.305 -25.885 -25.205 ;
      RECT -25.985 -25.065 -25.885 -24.965 ;
      RECT -25.985 -23.485 -25.885 -23.385 ;
      RECT -25.985 -23.245 -25.885 -23.145 ;
      RECT -25.985 -22.955 -25.885 -22.855 ;
      RECT -25.985 -18.725 -25.885 -18.625 ;
      RECT -25.985 -18.485 -25.885 -18.385 ;
      RECT -25.985 -17.145 -25.885 -17.045 ;
      RECT -25.985 -16.905 -25.885 -16.805 ;
      RECT -25.985 -12.675 -25.885 -12.575 ;
      RECT -25.985 -12.385 -25.885 -12.285 ;
      RECT -25.985 -12.145 -25.885 -12.045 ;
      RECT -25.985 -10.565 -25.885 -10.465 ;
      RECT -25.985 -10.325 -25.885 -10.225 ;
      RECT -25.985 -10.035 -25.885 -9.935 ;
      RECT -25.985 -5.805 -25.885 -5.705 ;
      RECT -25.985 -5.565 -25.885 -5.465 ;
      RECT -25.985 -4.225 -25.885 -4.125 ;
      RECT -25.985 -3.985 -25.885 -3.885 ;
      RECT -25.985 0.245 -25.885 0.345 ;
      RECT -25.985 0.535 -25.885 0.635 ;
      RECT -25.985 0.775 -25.885 0.875 ;
      RECT -26.825 -48.575 -26.725 -48.475 ;
      RECT -26.825 -38.735 -26.725 -38.635 ;
      RECT -26.825 -35.655 -26.725 -35.555 ;
      RECT -26.825 -25.815 -26.725 -25.715 ;
      RECT -26.825 -22.735 -26.725 -22.635 ;
      RECT -26.825 -12.895 -26.725 -12.795 ;
      RECT -26.825 -9.815 -26.725 -9.715 ;
      RECT -26.825 0.025 -26.725 0.125 ;
      RECT -26.865 2.235 -26.765 2.335 ;
      RECT -26.865 2.475 -26.765 2.575 ;
      RECT -26.865 4.895 -26.765 4.995 ;
      RECT -27.425 -48.135 -27.325 -48.035 ;
      RECT -27.425 -39.175 -27.325 -39.075 ;
      RECT -27.425 -35.215 -27.325 -35.115 ;
      RECT -27.425 -26.255 -27.325 -26.155 ;
      RECT -27.425 -22.295 -27.325 -22.195 ;
      RECT -27.425 -13.335 -27.325 -13.235 ;
      RECT -27.425 -9.375 -27.325 -9.275 ;
      RECT -27.425 -0.415 -27.325 -0.315 ;
      RECT -27.465 2.235 -27.365 2.335 ;
      RECT -27.465 2.475 -27.365 2.575 ;
      RECT -27.465 4.895 -27.365 4.995 ;
      RECT -28.025 -39.615 -27.925 -39.515 ;
      RECT -28.025 -26.695 -27.925 -26.595 ;
      RECT -28.025 -13.775 -27.925 -13.675 ;
      RECT -28.025 -0.855 -27.925 -0.755 ;
      RECT -28.065 2.235 -27.965 2.335 ;
      RECT -28.065 2.475 -27.965 2.575 ;
      RECT -28.065 4.895 -27.965 4.995 ;
      RECT -28.625 -34.555 -28.525 -34.455 ;
      RECT -28.625 -26.915 -28.525 -26.815 ;
      RECT -28.625 -8.715 -28.525 -8.615 ;
      RECT -28.625 -1.075 -28.525 -0.975 ;
      RECT -28.665 2.235 -28.565 2.335 ;
      RECT -28.665 2.475 -28.565 2.575 ;
      RECT -28.665 4.895 -28.565 4.995 ;
      RECT -29.225 -21.415 -29.125 -21.315 ;
      RECT -29.225 -14.215 -29.125 -14.115 ;
      RECT -29.225 -8.495 -29.125 -8.395 ;
      RECT -29.225 -1.295 -29.125 -1.195 ;
      RECT -29.265 2.235 -29.165 2.335 ;
      RECT -29.265 2.475 -29.165 2.575 ;
      RECT -29.265 4.895 -29.165 4.995 ;
    LAYER M2 ;
      RECT 36.545 -58.095 36.68 -57.595 ;
      RECT 36.545 -58.095 37.825 -57.99 ;
      RECT 37.725 -60.525 37.825 -57.99 ;
      RECT 36.21 -58.095 36.355 -57.595 ;
      RECT 35.705 -58.095 36.355 -57.99 ;
      RECT 35.705 -60.525 35.805 -57.99 ;
      RECT 34.675 -61.32 34.775 -55.535 ;
      RECT 34.315 -61.32 34.775 -61.22 ;
      RECT 34.315 -61.79 34.415 -61.22 ;
      RECT 33.965 -60.335 34.065 -58.875 ;
      RECT 33.925 -59.815 34.105 -59.715 ;
      RECT 31.745 -58.095 31.88 -57.595 ;
      RECT 31.745 -58.095 33.025 -57.99 ;
      RECT 32.925 -60.525 33.025 -57.99 ;
      RECT 31.41 -58.095 31.555 -57.595 ;
      RECT 30.905 -58.095 31.555 -57.99 ;
      RECT 30.905 -60.525 31.005 -57.99 ;
      RECT 29.875 -61.32 29.975 -55.535 ;
      RECT 29.515 -61.32 29.975 -61.22 ;
      RECT 29.515 -61.79 29.615 -61.22 ;
      RECT 29.165 -60.335 29.265 -58.875 ;
      RECT 29.125 -59.815 29.305 -59.715 ;
      RECT 26.945 -58.095 27.08 -57.595 ;
      RECT 26.945 -58.095 28.225 -57.99 ;
      RECT 28.125 -60.525 28.225 -57.99 ;
      RECT 26.61 -58.095 26.755 -57.595 ;
      RECT 26.105 -58.095 26.755 -57.99 ;
      RECT 26.105 -60.525 26.205 -57.99 ;
      RECT 25.075 -61.32 25.175 -55.535 ;
      RECT 24.715 -61.32 25.175 -61.22 ;
      RECT 24.715 -61.79 24.815 -61.22 ;
      RECT 24.365 -60.335 24.465 -58.875 ;
      RECT 24.325 -59.815 24.505 -59.715 ;
      RECT 22.145 -58.095 22.28 -57.595 ;
      RECT 22.145 -58.095 23.425 -57.99 ;
      RECT 23.325 -60.525 23.425 -57.99 ;
      RECT 21.81 -58.095 21.955 -57.595 ;
      RECT 21.305 -58.095 21.955 -57.99 ;
      RECT 21.305 -60.525 21.405 -57.99 ;
      RECT 20.275 -61.32 20.375 -55.535 ;
      RECT 19.915 -61.32 20.375 -61.22 ;
      RECT 19.915 -61.79 20.015 -61.22 ;
      RECT 19.565 -60.335 19.665 -58.875 ;
      RECT 19.525 -59.815 19.705 -59.715 ;
      RECT 17.345 -58.095 17.48 -57.595 ;
      RECT 17.345 -58.095 18.625 -57.99 ;
      RECT 18.525 -60.525 18.625 -57.99 ;
      RECT 17.01 -58.095 17.155 -57.595 ;
      RECT 16.505 -58.095 17.155 -57.99 ;
      RECT 16.505 -60.525 16.605 -57.99 ;
      RECT 15.475 -61.32 15.575 -55.535 ;
      RECT 15.115 -61.32 15.575 -61.22 ;
      RECT 15.115 -61.79 15.215 -61.22 ;
      RECT 14.765 -60.335 14.865 -58.875 ;
      RECT 14.725 -59.815 14.905 -59.715 ;
      RECT 12.545 -58.095 12.68 -57.595 ;
      RECT 12.545 -58.095 13.825 -57.99 ;
      RECT 13.725 -60.525 13.825 -57.99 ;
      RECT 12.21 -58.095 12.355 -57.595 ;
      RECT 11.705 -58.095 12.355 -57.99 ;
      RECT 11.705 -60.525 11.805 -57.99 ;
      RECT 10.675 -61.32 10.775 -55.535 ;
      RECT 10.315 -61.32 10.775 -61.22 ;
      RECT 10.315 -61.79 10.415 -61.22 ;
      RECT 9.965 -60.335 10.065 -58.875 ;
      RECT 9.925 -59.815 10.105 -59.715 ;
      RECT 7.745 -58.095 7.88 -57.595 ;
      RECT 7.745 -58.095 9.025 -57.99 ;
      RECT 8.925 -60.525 9.025 -57.99 ;
      RECT 7.41 -58.095 7.555 -57.595 ;
      RECT 6.905 -58.095 7.555 -57.99 ;
      RECT 6.905 -60.525 7.005 -57.99 ;
      RECT 5.875 -61.32 5.975 -55.535 ;
      RECT 5.515 -61.32 5.975 -61.22 ;
      RECT 5.515 -61.79 5.615 -61.22 ;
      RECT 5.165 -60.335 5.265 -58.875 ;
      RECT 5.125 -59.815 5.305 -59.715 ;
      RECT 2.945 -58.095 3.08 -57.595 ;
      RECT 2.945 -58.095 4.225 -57.99 ;
      RECT 4.125 -60.525 4.225 -57.99 ;
      RECT 2.61 -58.095 2.755 -57.595 ;
      RECT 2.105 -58.095 2.755 -57.99 ;
      RECT 2.105 -60.525 2.205 -57.99 ;
      RECT 1.075 -61.32 1.175 -55.535 ;
      RECT 0.715 -61.32 1.175 -61.22 ;
      RECT 0.715 -61.79 0.815 -61.22 ;
      RECT 0.365 -60.335 0.465 -58.875 ;
      RECT 0.325 -59.815 0.505 -59.715 ;
      RECT -11.265 -55.495 -11.085 -51.035 ;
      RECT -11.265 -58.955 -11.165 -51.035 ;
      RECT -11.865 -55.495 -11.685 -51.035 ;
      RECT -11.865 -58.955 -11.765 -51.035 ;
      RECT -26.865 -49.035 -26.765 5.065 ;
      RECT -26.865 -49.035 -26.685 0.645 ;
      RECT -27.465 -49.035 -27.365 5.065 ;
      RECT -27.465 -49.035 -27.285 0.645 ;
      RECT -28.065 -49.035 -27.965 5.065 ;
      RECT -28.065 -49.035 -27.885 0.645 ;
      RECT -28.665 -49.035 -28.565 5.065 ;
      RECT -28.665 -49.035 -28.485 0.645 ;
      RECT -29.265 -49.035 -29.165 5.065 ;
      RECT -29.265 -49.035 -29.085 0.645 ;
      RECT 38.275 -57.285 38.375 -52.305 ;
      RECT 38.015 -53.265 38.115 3.135 ;
      RECT 37.585 -53.265 37.685 3.135 ;
      RECT 37.325 -57.005 37.425 -52.305 ;
      RECT 37.135 -60.305 37.235 -58.69 ;
      RECT 37.075 -57.285 37.175 -52.305 ;
      RECT 36.835 -57.51 36.935 -56.825 ;
      RECT 36.815 -53.265 36.915 3.135 ;
      RECT 36.385 -53.265 36.485 3.135 ;
      RECT 36.125 -57.005 36.225 -52.305 ;
      RECT 35.875 -57.285 35.975 -55.535 ;
      RECT 35.615 -56.495 35.715 3.135 ;
      RECT 35.185 -56.495 35.285 3.135 ;
      RECT 35.115 -60.305 35.215 -58.705 ;
      RECT 34.925 -57.005 35.025 -55.535 ;
      RECT 34.415 -56.495 34.515 3.135 ;
      RECT 33.985 -56.495 34.085 3.135 ;
      RECT 33.725 -61.79 33.825 -55.535 ;
      RECT 33.475 -57.285 33.575 -52.305 ;
      RECT 33.215 -53.265 33.315 3.135 ;
      RECT 32.785 -53.265 32.885 3.135 ;
      RECT 32.525 -57.005 32.625 -52.305 ;
      RECT 32.335 -60.305 32.435 -58.69 ;
      RECT 32.275 -57.285 32.375 -52.305 ;
      RECT 32.035 -57.51 32.135 -56.825 ;
      RECT 32.015 -53.265 32.115 3.135 ;
      RECT 31.585 -53.265 31.685 3.135 ;
      RECT 31.325 -57.005 31.425 -52.305 ;
      RECT 31.075 -57.285 31.175 -55.535 ;
      RECT 30.815 -56.495 30.915 3.135 ;
      RECT 30.385 -56.495 30.485 3.135 ;
      RECT 30.315 -60.305 30.415 -58.705 ;
      RECT 30.125 -57.005 30.225 -55.535 ;
      RECT 29.615 -56.495 29.715 3.135 ;
      RECT 29.185 -56.495 29.285 3.135 ;
      RECT 28.925 -61.79 29.025 -55.535 ;
      RECT 28.675 -57.285 28.775 -52.305 ;
      RECT 28.415 -53.265 28.515 3.135 ;
      RECT 27.985 -53.265 28.085 3.135 ;
      RECT 27.725 -57.005 27.825 -52.305 ;
      RECT 27.535 -60.305 27.635 -58.69 ;
      RECT 27.475 -57.285 27.575 -52.305 ;
      RECT 27.235 -57.51 27.335 -56.825 ;
      RECT 27.215 -53.265 27.315 3.135 ;
      RECT 26.785 -53.265 26.885 3.135 ;
      RECT 26.525 -57.005 26.625 -52.305 ;
      RECT 26.275 -57.285 26.375 -55.535 ;
      RECT 26.015 -56.495 26.115 3.135 ;
      RECT 25.585 -56.495 25.685 3.135 ;
      RECT 25.515 -60.305 25.615 -58.705 ;
      RECT 25.325 -57.005 25.425 -55.535 ;
      RECT 24.815 -56.495 24.915 3.135 ;
      RECT 24.385 -56.495 24.485 3.135 ;
      RECT 24.125 -61.79 24.225 -55.535 ;
      RECT 23.875 -57.285 23.975 -52.305 ;
      RECT 23.615 -53.265 23.715 3.135 ;
      RECT 23.185 -53.265 23.285 3.135 ;
      RECT 22.925 -57.005 23.025 -52.305 ;
      RECT 22.735 -60.305 22.835 -58.69 ;
      RECT 22.675 -57.285 22.775 -52.305 ;
      RECT 22.435 -57.51 22.535 -56.825 ;
      RECT 22.415 -53.265 22.515 3.135 ;
      RECT 21.985 -53.265 22.085 3.135 ;
      RECT 21.725 -57.005 21.825 -52.305 ;
      RECT 21.475 -57.285 21.575 -55.535 ;
      RECT 21.215 -56.495 21.315 3.135 ;
      RECT 20.785 -56.495 20.885 3.135 ;
      RECT 20.715 -60.305 20.815 -58.705 ;
      RECT 20.525 -57.005 20.625 -55.535 ;
      RECT 20.015 -56.495 20.115 3.135 ;
      RECT 19.585 -56.495 19.685 3.135 ;
      RECT 19.325 -61.79 19.425 -55.535 ;
      RECT 19.075 -57.285 19.175 -52.305 ;
      RECT 18.815 -53.265 18.915 3.135 ;
      RECT 18.385 -53.265 18.485 3.135 ;
      RECT 18.125 -57.005 18.225 -52.305 ;
      RECT 17.935 -60.305 18.035 -58.69 ;
      RECT 17.875 -57.285 17.975 -52.305 ;
      RECT 17.635 -57.51 17.735 -56.825 ;
      RECT 17.615 -53.265 17.715 3.135 ;
      RECT 17.185 -53.265 17.285 3.135 ;
      RECT 16.925 -57.005 17.025 -52.305 ;
      RECT 16.675 -57.285 16.775 -55.535 ;
      RECT 16.415 -56.495 16.515 3.135 ;
      RECT 15.985 -56.495 16.085 3.135 ;
      RECT 15.915 -60.305 16.015 -58.705 ;
      RECT 15.725 -57.005 15.825 -55.535 ;
      RECT 15.215 -56.495 15.315 3.135 ;
      RECT 14.785 -56.495 14.885 3.135 ;
      RECT 14.525 -61.79 14.625 -55.535 ;
      RECT 14.275 -57.285 14.375 -52.305 ;
      RECT 14.015 -53.265 14.115 3.135 ;
      RECT 13.585 -53.265 13.685 3.135 ;
      RECT 13.325 -57.005 13.425 -52.305 ;
      RECT 13.135 -60.305 13.235 -58.69 ;
      RECT 13.075 -57.285 13.175 -52.305 ;
      RECT 12.835 -57.51 12.935 -56.825 ;
      RECT 12.815 -53.265 12.915 3.135 ;
      RECT 12.385 -53.265 12.485 3.135 ;
      RECT 12.125 -57.005 12.225 -52.305 ;
      RECT 11.875 -57.285 11.975 -55.535 ;
      RECT 11.615 -56.495 11.715 3.135 ;
      RECT 11.185 -56.495 11.285 3.135 ;
      RECT 11.115 -60.305 11.215 -58.705 ;
      RECT 10.925 -57.005 11.025 -55.535 ;
      RECT 10.415 -56.495 10.515 3.135 ;
      RECT 9.985 -56.495 10.085 3.135 ;
      RECT 9.725 -61.79 9.825 -55.535 ;
      RECT 9.475 -57.285 9.575 -52.305 ;
      RECT 9.215 -53.265 9.315 3.135 ;
      RECT 8.785 -53.265 8.885 3.135 ;
      RECT 8.525 -57.005 8.625 -52.305 ;
      RECT 8.335 -60.305 8.435 -58.69 ;
      RECT 8.275 -57.285 8.375 -52.305 ;
      RECT 8.035 -57.51 8.135 -56.825 ;
      RECT 8.015 -53.265 8.115 3.135 ;
      RECT 7.585 -53.265 7.685 3.135 ;
      RECT 7.325 -57.005 7.425 -52.305 ;
      RECT 7.075 -57.285 7.175 -55.535 ;
      RECT 6.815 -56.495 6.915 3.135 ;
      RECT 6.385 -56.495 6.485 3.135 ;
      RECT 6.315 -60.305 6.415 -58.705 ;
      RECT 6.125 -57.005 6.225 -55.535 ;
      RECT 5.615 -56.495 5.715 3.135 ;
      RECT 5.185 -56.495 5.285 3.135 ;
      RECT 4.925 -61.79 5.025 -55.535 ;
      RECT 4.675 -57.285 4.775 -52.305 ;
      RECT 4.415 -53.265 4.515 3.135 ;
      RECT 3.985 -53.265 4.085 3.135 ;
      RECT 3.725 -57.005 3.825 -52.305 ;
      RECT 3.535 -60.305 3.635 -58.69 ;
      RECT 3.475 -57.285 3.575 -52.305 ;
      RECT 3.235 -57.51 3.335 -56.825 ;
      RECT 3.215 -53.265 3.315 3.135 ;
      RECT 2.785 -53.265 2.885 3.135 ;
      RECT 2.525 -57.005 2.625 -52.305 ;
      RECT 2.275 -57.285 2.375 -55.535 ;
      RECT 2.015 -56.495 2.115 3.135 ;
      RECT 1.585 -56.495 1.685 3.135 ;
      RECT 1.515 -60.305 1.615 -58.705 ;
      RECT 1.325 -57.005 1.425 -55.535 ;
      RECT 0.815 -56.495 0.915 3.135 ;
      RECT 0.385 -56.495 0.485 3.135 ;
      RECT 0.125 -61.79 0.225 -55.535 ;
      RECT -0.385 1.895 -0.285 4.275 ;
      RECT -0.765 -55.975 -0.665 -50.615 ;
      RECT -0.765 -49.515 -0.665 -44.155 ;
      RECT -0.765 -43.055 -0.665 -37.695 ;
      RECT -0.765 -36.595 -0.665 -31.235 ;
      RECT -0.765 -30.135 -0.665 -24.775 ;
      RECT -0.765 -23.675 -0.665 -18.315 ;
      RECT -0.765 -17.215 -0.665 -11.855 ;
      RECT -0.765 -10.755 -0.665 -5.395 ;
      RECT -0.765 -4.295 -0.665 1.065 ;
      RECT -1.285 -55.975 -1.185 -50.615 ;
      RECT -1.285 -49.515 -1.185 -44.155 ;
      RECT -1.285 -43.055 -1.185 -37.695 ;
      RECT -1.285 -36.595 -1.185 -31.235 ;
      RECT -1.285 -30.135 -1.185 -24.775 ;
      RECT -1.285 -23.675 -1.185 -18.315 ;
      RECT -1.285 -17.215 -1.185 -11.855 ;
      RECT -1.285 -10.755 -1.185 -5.395 ;
      RECT -1.285 -4.295 -1.185 1.065 ;
      RECT -1.805 -51.77 -1.705 -50.615 ;
      RECT -1.805 -49.515 -1.705 -48.36 ;
      RECT -1.805 -38.85 -1.705 -37.695 ;
      RECT -1.805 -36.595 -1.705 -35.44 ;
      RECT -1.805 -25.93 -1.705 -24.775 ;
      RECT -1.805 -23.675 -1.705 -22.52 ;
      RECT -1.805 -13.01 -1.705 -11.855 ;
      RECT -1.805 -10.755 -1.705 -9.6 ;
      RECT -1.805 -0.09 -1.705 1.065 ;
      RECT -2.065 -55.975 -1.965 -50.615 ;
      RECT -2.065 -49.515 -1.965 -44.155 ;
      RECT -2.065 -43.055 -1.965 -37.695 ;
      RECT -2.065 -36.595 -1.965 -31.235 ;
      RECT -2.065 -30.135 -1.965 -24.775 ;
      RECT -2.065 -23.675 -1.965 -18.315 ;
      RECT -2.065 -17.215 -1.965 -11.855 ;
      RECT -2.065 -10.755 -1.965 -5.395 ;
      RECT -2.065 -4.295 -1.965 1.065 ;
      RECT -2.585 -55.975 -2.485 -50.615 ;
      RECT -2.585 -49.515 -2.485 -44.155 ;
      RECT -2.585 -43.055 -2.485 -37.695 ;
      RECT -2.585 -36.595 -2.485 -31.235 ;
      RECT -2.585 -30.135 -2.485 -24.775 ;
      RECT -2.585 -23.675 -2.485 -18.315 ;
      RECT -2.585 -17.215 -2.485 -11.855 ;
      RECT -2.585 -10.755 -2.485 -5.395 ;
      RECT -2.585 -4.295 -2.485 1.065 ;
      RECT -3.105 -51.77 -3.005 -50.615 ;
      RECT -3.105 -49.515 -3.005 -48.36 ;
      RECT -3.105 -38.85 -3.005 -37.695 ;
      RECT -3.105 -36.595 -3.005 -35.44 ;
      RECT -3.105 -25.93 -3.005 -24.775 ;
      RECT -3.105 -23.675 -3.005 -22.52 ;
      RECT -3.105 -13.01 -3.005 -11.855 ;
      RECT -3.105 -10.755 -3.005 -9.6 ;
      RECT -3.105 -0.09 -3.005 1.065 ;
      RECT -3.365 -55.975 -3.265 -50.615 ;
      RECT -3.365 -49.515 -3.265 -44.155 ;
      RECT -3.365 -43.055 -3.265 -37.695 ;
      RECT -3.365 -36.595 -3.265 -31.235 ;
      RECT -3.365 -30.135 -3.265 -24.775 ;
      RECT -3.365 -23.675 -3.265 -18.315 ;
      RECT -3.365 -17.215 -3.265 -11.855 ;
      RECT -3.365 -10.755 -3.265 -5.395 ;
      RECT -3.365 -4.295 -3.265 1.065 ;
      RECT -3.885 -55.975 -3.785 -50.615 ;
      RECT -3.885 -49.515 -3.785 -44.155 ;
      RECT -3.885 -43.055 -3.785 -37.695 ;
      RECT -3.885 -36.595 -3.785 -31.235 ;
      RECT -3.885 -30.135 -3.785 -24.775 ;
      RECT -3.885 -23.675 -3.785 -18.315 ;
      RECT -3.885 -17.215 -3.785 -11.855 ;
      RECT -3.885 -10.755 -3.785 -5.395 ;
      RECT -3.885 -4.295 -3.785 1.065 ;
      RECT -4.405 -51.77 -4.305 -50.615 ;
      RECT -4.405 -49.515 -4.305 -48.36 ;
      RECT -4.405 -38.85 -4.305 -37.695 ;
      RECT -4.405 -36.595 -4.305 -35.44 ;
      RECT -4.405 -25.93 -4.305 -24.775 ;
      RECT -4.405 -23.675 -4.305 -22.52 ;
      RECT -4.405 -13.01 -4.305 -11.855 ;
      RECT -4.405 -10.755 -4.305 -9.6 ;
      RECT -4.405 -0.09 -4.305 1.065 ;
      RECT -4.665 -55.975 -4.565 -50.615 ;
      RECT -4.665 -49.515 -4.565 -44.155 ;
      RECT -4.665 -43.055 -4.565 -37.695 ;
      RECT -4.665 -36.595 -4.565 -31.235 ;
      RECT -4.665 -30.135 -4.565 -24.775 ;
      RECT -4.665 -23.675 -4.565 -18.315 ;
      RECT -4.665 -17.215 -4.565 -11.855 ;
      RECT -4.665 -10.755 -4.565 -5.395 ;
      RECT -4.665 -4.295 -4.565 1.065 ;
      RECT -4.925 -59.535 -4.825 4.275 ;
      RECT -5.185 -55.975 -5.085 -50.615 ;
      RECT -5.185 -49.515 -5.085 -44.155 ;
      RECT -5.185 -43.055 -5.085 -37.695 ;
      RECT -5.185 -36.595 -5.085 -31.235 ;
      RECT -5.185 -30.135 -5.085 -24.775 ;
      RECT -5.185 -23.675 -5.085 -18.315 ;
      RECT -5.185 -17.215 -5.085 -11.855 ;
      RECT -5.185 -10.755 -5.085 -5.395 ;
      RECT -5.185 -4.295 -5.085 1.065 ;
      RECT -5.705 -51.77 -5.605 -50.615 ;
      RECT -5.705 -49.515 -5.605 -48.36 ;
      RECT -5.705 -38.85 -5.605 -37.695 ;
      RECT -5.705 -36.595 -5.605 -35.44 ;
      RECT -5.705 -25.93 -5.605 -24.775 ;
      RECT -5.705 -23.675 -5.605 -22.52 ;
      RECT -5.705 -13.01 -5.605 -11.855 ;
      RECT -5.705 -10.755 -5.605 -9.6 ;
      RECT -5.705 -0.09 -5.605 1.065 ;
      RECT -5.965 -55.975 -5.865 -50.615 ;
      RECT -5.965 -49.515 -5.865 -44.155 ;
      RECT -5.965 -43.055 -5.865 -37.695 ;
      RECT -5.965 -36.595 -5.865 -31.235 ;
      RECT -5.965 -30.135 -5.865 -24.775 ;
      RECT -5.965 -23.675 -5.865 -18.315 ;
      RECT -5.965 -17.215 -5.865 -11.855 ;
      RECT -5.965 -10.755 -5.865 -5.395 ;
      RECT -5.965 -4.295 -5.865 1.065 ;
      RECT -6.485 -55.975 -6.385 -50.615 ;
      RECT -6.485 -49.515 -6.385 -44.155 ;
      RECT -6.485 -43.055 -6.385 -37.695 ;
      RECT -6.485 -36.595 -6.385 -31.235 ;
      RECT -6.485 -30.135 -6.385 -24.775 ;
      RECT -6.485 -23.675 -6.385 -18.315 ;
      RECT -6.485 -17.215 -6.385 -11.855 ;
      RECT -6.485 -10.755 -6.385 -5.395 ;
      RECT -6.485 -4.295 -6.385 1.065 ;
      RECT -7.265 -55.975 -7.165 -50.615 ;
      RECT -7.265 -49.515 -7.165 -44.155 ;
      RECT -7.265 -43.055 -7.165 -37.695 ;
      RECT -7.265 -36.595 -7.165 -31.235 ;
      RECT -7.265 -30.135 -7.165 -24.775 ;
      RECT -7.265 -23.675 -7.165 -18.315 ;
      RECT -7.265 -17.215 -7.165 -11.855 ;
      RECT -7.265 -10.755 -7.165 -5.395 ;
      RECT -7.265 -4.295 -7.165 1.065 ;
      RECT -7.785 -55.975 -7.685 -50.615 ;
      RECT -7.785 -49.515 -7.685 -44.155 ;
      RECT -7.785 -43.055 -7.685 -37.695 ;
      RECT -7.785 -36.595 -7.685 -31.235 ;
      RECT -7.785 -30.135 -7.685 -24.775 ;
      RECT -7.785 -23.675 -7.685 -18.315 ;
      RECT -7.785 -17.215 -7.685 -11.855 ;
      RECT -7.785 -10.755 -7.685 -5.395 ;
      RECT -7.785 -4.295 -7.685 1.065 ;
      RECT -8.565 -55.975 -8.465 -50.615 ;
      RECT -8.565 -49.515 -8.465 -44.155 ;
      RECT -8.565 -43.055 -8.465 -37.695 ;
      RECT -8.565 -36.595 -8.465 -31.235 ;
      RECT -8.565 -30.135 -8.465 -24.775 ;
      RECT -8.565 -23.675 -8.465 -18.315 ;
      RECT -8.565 -17.215 -8.465 -11.855 ;
      RECT -8.565 -10.755 -8.465 -5.395 ;
      RECT -8.565 -4.295 -8.465 1.065 ;
      RECT -9.085 -55.975 -8.985 -50.615 ;
      RECT -9.085 -49.515 -8.985 -44.155 ;
      RECT -9.085 -43.055 -8.985 -37.695 ;
      RECT -9.085 -36.595 -8.985 -31.235 ;
      RECT -9.085 -30.135 -8.985 -24.775 ;
      RECT -9.085 -23.675 -8.985 -18.315 ;
      RECT -9.085 -17.215 -8.985 -11.855 ;
      RECT -9.085 -10.755 -8.985 -5.395 ;
      RECT -9.085 -4.295 -8.985 1.065 ;
      RECT -9.865 -55.975 -9.765 -50.615 ;
      RECT -9.865 -49.515 -9.765 -44.155 ;
      RECT -9.865 -43.055 -9.765 -37.695 ;
      RECT -9.865 -36.595 -9.765 -31.235 ;
      RECT -9.865 -30.135 -9.765 -24.775 ;
      RECT -9.865 -23.675 -9.765 -18.315 ;
      RECT -9.865 -17.215 -9.765 -11.855 ;
      RECT -9.865 -10.755 -9.765 -5.395 ;
      RECT -9.865 -4.295 -9.765 1.065 ;
      RECT -10.385 -55.975 -10.285 -50.615 ;
      RECT -10.385 -49.515 -10.285 -44.155 ;
      RECT -10.385 -43.055 -10.285 -37.695 ;
      RECT -10.385 -36.595 -10.285 -31.235 ;
      RECT -10.385 -30.135 -10.285 -24.775 ;
      RECT -10.385 -23.675 -10.285 -18.315 ;
      RECT -10.385 -17.215 -10.285 -11.855 ;
      RECT -10.385 -10.755 -10.285 -5.395 ;
      RECT -10.385 -4.295 -10.285 1.065 ;
      RECT -11.165 -49.515 -11.065 -44.155 ;
      RECT -11.165 -43.055 -11.065 -37.695 ;
      RECT -11.165 -36.595 -11.065 -31.235 ;
      RECT -11.165 -30.135 -11.065 -24.775 ;
      RECT -11.165 -23.675 -11.065 -18.315 ;
      RECT -11.165 -17.215 -11.065 -11.855 ;
      RECT -11.165 -10.755 -11.065 -5.395 ;
      RECT -11.165 -4.295 -11.065 1.065 ;
      RECT -11.685 -49.515 -11.585 -44.155 ;
      RECT -11.685 -43.055 -11.585 -37.695 ;
      RECT -11.685 -36.595 -11.585 -31.235 ;
      RECT -11.685 -30.135 -11.585 -24.775 ;
      RECT -11.685 -23.675 -11.585 -18.315 ;
      RECT -11.685 -17.215 -11.585 -11.855 ;
      RECT -11.685 -10.755 -11.585 -5.395 ;
      RECT -11.685 -4.295 -11.585 1.065 ;
      RECT -12.465 -49.515 -12.365 -44.155 ;
      RECT -12.465 -43.055 -12.365 -37.695 ;
      RECT -12.465 -36.595 -12.365 -31.235 ;
      RECT -12.465 -30.135 -12.365 -24.775 ;
      RECT -12.465 -23.675 -12.365 -18.315 ;
      RECT -12.465 -17.215 -12.365 -11.855 ;
      RECT -12.465 -10.755 -12.365 -5.395 ;
      RECT -12.465 -4.295 -12.365 1.065 ;
      RECT -12.985 -49.515 -12.885 -44.155 ;
      RECT -12.985 -43.055 -12.885 -37.695 ;
      RECT -12.985 -36.595 -12.885 -31.235 ;
      RECT -12.985 -30.135 -12.885 -24.775 ;
      RECT -12.985 -23.675 -12.885 -18.315 ;
      RECT -12.985 -17.215 -12.885 -11.855 ;
      RECT -12.985 -10.755 -12.885 -5.395 ;
      RECT -12.985 -4.295 -12.885 1.065 ;
      RECT -13.765 -49.515 -13.665 -44.155 ;
      RECT -13.765 -43.055 -13.665 -37.695 ;
      RECT -13.765 -36.595 -13.665 -31.235 ;
      RECT -13.765 -30.135 -13.665 -24.775 ;
      RECT -13.765 -23.675 -13.665 -18.315 ;
      RECT -13.765 -17.215 -13.665 -11.855 ;
      RECT -13.765 -10.755 -13.665 -5.395 ;
      RECT -13.765 -4.295 -13.665 1.065 ;
      RECT -14.285 -49.515 -14.185 -44.155 ;
      RECT -14.285 -43.055 -14.185 -37.695 ;
      RECT -14.285 -36.595 -14.185 -31.235 ;
      RECT -14.285 -30.135 -14.185 -24.775 ;
      RECT -14.285 -23.675 -14.185 -18.315 ;
      RECT -14.285 -17.215 -14.185 -11.855 ;
      RECT -14.285 -10.755 -14.185 -5.395 ;
      RECT -14.285 -4.295 -14.185 1.065 ;
      RECT -15.065 -49.515 -14.965 -44.155 ;
      RECT -15.065 -43.055 -14.965 -37.695 ;
      RECT -15.065 -36.595 -14.965 -31.235 ;
      RECT -15.065 -30.135 -14.965 -24.775 ;
      RECT -15.065 -23.675 -14.965 -18.315 ;
      RECT -15.065 -17.215 -14.965 -11.855 ;
      RECT -15.065 -10.755 -14.965 -5.395 ;
      RECT -15.065 -4.295 -14.965 1.065 ;
      RECT -15.585 -49.515 -15.485 -44.155 ;
      RECT -15.585 -43.055 -15.485 -37.695 ;
      RECT -15.585 -36.595 -15.485 -31.235 ;
      RECT -15.585 -30.135 -15.485 -24.775 ;
      RECT -15.585 -23.675 -15.485 -18.315 ;
      RECT -15.585 -17.215 -15.485 -11.855 ;
      RECT -15.585 -10.755 -15.485 -5.395 ;
      RECT -15.585 -4.295 -15.485 1.065 ;
      RECT -16.365 -49.515 -16.265 -44.155 ;
      RECT -16.365 -43.055 -16.265 -37.695 ;
      RECT -16.365 -36.595 -16.265 -31.235 ;
      RECT -16.365 -30.135 -16.265 -24.775 ;
      RECT -16.365 -23.675 -16.265 -18.315 ;
      RECT -16.365 -17.215 -16.265 -11.855 ;
      RECT -16.365 -10.755 -16.265 -5.395 ;
      RECT -16.365 -4.295 -16.265 1.065 ;
      RECT -16.885 -49.515 -16.785 -44.155 ;
      RECT -16.885 -43.055 -16.785 -37.695 ;
      RECT -16.885 -36.595 -16.785 -31.235 ;
      RECT -16.885 -30.135 -16.785 -24.775 ;
      RECT -16.885 -23.675 -16.785 -18.315 ;
      RECT -16.885 -17.215 -16.785 -11.855 ;
      RECT -16.885 -10.755 -16.785 -5.395 ;
      RECT -16.885 -4.295 -16.785 1.065 ;
      RECT -17.665 -49.515 -17.565 -44.155 ;
      RECT -17.665 -43.055 -17.565 -37.695 ;
      RECT -17.665 -36.595 -17.565 -31.235 ;
      RECT -17.665 -30.135 -17.565 -24.775 ;
      RECT -17.665 -23.675 -17.565 -18.315 ;
      RECT -17.665 -17.215 -17.565 -11.855 ;
      RECT -17.665 -10.755 -17.565 -5.395 ;
      RECT -17.665 -4.295 -17.565 1.065 ;
      RECT -18.185 -49.515 -18.085 -44.155 ;
      RECT -18.185 -43.055 -18.085 -37.695 ;
      RECT -18.185 -36.595 -18.085 -31.235 ;
      RECT -18.185 -30.135 -18.085 -24.775 ;
      RECT -18.185 -23.675 -18.085 -18.315 ;
      RECT -18.185 -17.215 -18.085 -11.855 ;
      RECT -18.185 -10.755 -18.085 -5.395 ;
      RECT -18.185 -4.295 -18.085 1.065 ;
      RECT -18.965 -49.515 -18.865 -44.155 ;
      RECT -18.965 -43.055 -18.865 -37.695 ;
      RECT -18.965 -36.595 -18.865 -31.235 ;
      RECT -18.965 -30.135 -18.865 -24.775 ;
      RECT -18.965 -23.675 -18.865 -18.315 ;
      RECT -18.965 -17.215 -18.865 -11.855 ;
      RECT -18.965 -10.755 -18.865 -5.395 ;
      RECT -18.965 -4.295 -18.865 1.065 ;
      RECT -19.485 -49.515 -19.385 -44.155 ;
      RECT -19.485 -43.055 -19.385 -37.695 ;
      RECT -19.485 -36.595 -19.385 -31.235 ;
      RECT -19.485 -30.135 -19.385 -24.775 ;
      RECT -19.485 -23.675 -19.385 -18.315 ;
      RECT -19.485 -17.215 -19.385 -11.855 ;
      RECT -19.485 -10.755 -19.385 -5.395 ;
      RECT -19.485 -4.295 -19.385 1.065 ;
      RECT -20.265 -49.515 -20.165 -44.155 ;
      RECT -20.265 -43.055 -20.165 -37.695 ;
      RECT -20.265 -36.595 -20.165 -31.235 ;
      RECT -20.265 -30.135 -20.165 -24.775 ;
      RECT -20.265 -23.675 -20.165 -18.315 ;
      RECT -20.265 -17.215 -20.165 -11.855 ;
      RECT -20.265 -10.755 -20.165 -5.395 ;
      RECT -20.265 -4.295 -20.165 1.065 ;
      RECT -20.785 -49.515 -20.685 -44.155 ;
      RECT -20.785 -43.055 -20.685 -37.695 ;
      RECT -20.785 -36.595 -20.685 -31.235 ;
      RECT -20.785 -30.135 -20.685 -24.775 ;
      RECT -20.785 -23.675 -20.685 -18.315 ;
      RECT -20.785 -17.215 -20.685 -11.855 ;
      RECT -20.785 -10.755 -20.685 -5.395 ;
      RECT -20.785 -4.295 -20.685 1.065 ;
      RECT -21.565 -49.515 -21.465 -44.155 ;
      RECT -21.565 -43.055 -21.465 -37.695 ;
      RECT -21.565 -36.595 -21.465 -31.235 ;
      RECT -21.565 -30.135 -21.465 -24.775 ;
      RECT -21.565 -23.675 -21.465 -18.315 ;
      RECT -21.565 -17.215 -21.465 -11.855 ;
      RECT -21.565 -10.755 -21.465 -5.395 ;
      RECT -21.565 -4.295 -21.465 1.065 ;
      RECT -22.085 -49.515 -21.985 -44.155 ;
      RECT -22.085 -43.055 -21.985 -37.695 ;
      RECT -22.085 -36.595 -21.985 -31.235 ;
      RECT -22.085 -30.135 -21.985 -24.775 ;
      RECT -22.085 -23.675 -21.985 -18.315 ;
      RECT -22.085 -17.215 -21.985 -11.855 ;
      RECT -22.085 -10.755 -21.985 -5.395 ;
      RECT -22.085 -4.295 -21.985 1.065 ;
      RECT -22.865 -49.515 -22.765 -44.155 ;
      RECT -22.865 -43.055 -22.765 -37.695 ;
      RECT -22.865 -36.595 -22.765 -31.235 ;
      RECT -22.865 -30.135 -22.765 -24.775 ;
      RECT -22.865 -23.675 -22.765 -18.315 ;
      RECT -22.865 -17.215 -22.765 -11.855 ;
      RECT -22.865 -10.755 -22.765 -5.395 ;
      RECT -22.865 -4.295 -22.765 1.065 ;
      RECT -23.385 -49.515 -23.285 -44.155 ;
      RECT -23.385 -43.055 -23.285 -37.695 ;
      RECT -23.385 -36.595 -23.285 -31.235 ;
      RECT -23.385 -30.135 -23.285 -24.775 ;
      RECT -23.385 -23.675 -23.285 -18.315 ;
      RECT -23.385 -17.215 -23.285 -11.855 ;
      RECT -23.385 -10.755 -23.285 -5.395 ;
      RECT -23.385 -4.295 -23.285 1.065 ;
      RECT -24.165 -49.515 -24.065 -44.155 ;
      RECT -24.165 -43.055 -24.065 -37.695 ;
      RECT -24.165 -36.595 -24.065 -31.235 ;
      RECT -24.165 -30.135 -24.065 -24.775 ;
      RECT -24.165 -23.675 -24.065 -18.315 ;
      RECT -24.165 -17.215 -24.065 -11.855 ;
      RECT -24.165 -10.755 -24.065 -5.395 ;
      RECT -24.165 -4.295 -24.065 1.065 ;
      RECT -24.685 -49.515 -24.585 -44.155 ;
      RECT -24.685 -43.055 -24.585 -37.695 ;
      RECT -24.685 -36.595 -24.585 -31.235 ;
      RECT -24.685 -30.135 -24.585 -24.775 ;
      RECT -24.685 -23.675 -24.585 -18.315 ;
      RECT -24.685 -17.215 -24.585 -11.855 ;
      RECT -24.685 -10.755 -24.585 -5.395 ;
      RECT -24.685 -4.295 -24.585 1.065 ;
      RECT -25.465 -49.515 -25.365 -44.155 ;
      RECT -25.465 -43.055 -25.365 -37.695 ;
      RECT -25.465 -36.595 -25.365 -31.235 ;
      RECT -25.465 -30.135 -25.365 -24.775 ;
      RECT -25.465 -23.675 -25.365 -18.315 ;
      RECT -25.465 -17.215 -25.365 -11.855 ;
      RECT -25.465 -10.755 -25.365 -5.395 ;
      RECT -25.465 -4.295 -25.365 1.065 ;
      RECT -25.985 -49.515 -25.885 -44.155 ;
      RECT -25.985 -43.055 -25.885 -37.695 ;
      RECT -25.985 -36.595 -25.885 -31.235 ;
      RECT -25.985 -30.135 -25.885 -24.775 ;
      RECT -25.985 -23.675 -25.885 -18.315 ;
      RECT -25.985 -17.215 -25.885 -11.855 ;
      RECT -25.985 -10.755 -25.885 -5.395 ;
      RECT -25.985 -4.295 -25.885 1.065 ;
  END
END sram_compiled_array

END LIBRARY
